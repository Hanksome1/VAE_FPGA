`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/06/13 22:33:04
// Design Name: 
// Module Name: decoder4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module decoder4 #(
    parameter output_number=10, 
    parameter input_number=200, 
    parameter width=11)(
    input clk, 
    input rst_n,
    input signed[width-1:0]input_node[0:input_number-1], 
    input enable, 
    output signed[width-1:0]output_node[0:output_number-1], 
    output finish
    );
wire signed [width-1:0] internode [0:output_number-1];
localparam signed [width-1:0] bias [0:output_number-1]= '{-12,-5,0,-1,-9,-5,-5,-7,-17,0,-3,5,-5,1,-6,-7,-9,3,-4,-12,-14,-15,-7,-13,1,0,5,-3,2,0,-5,0,-2,-1,-7,-14,7,11,0,6,-4,-5,-20,-16,-13,-5,15,22,21,33,26,29,7,0,-6,-14,-9,-25,0,14,24,15,16,17,6,16,11,-2,-11,-2,-4,-4,8,18,13,-13,1,-5,-17,6,-1,2,-22,-21,-10,-7,-1,11,-12,0,12,1,18,17,-5,-18,-10,-11,-8,-22,-11,16,16,31,27,22,37,12,-7,-8,1,-15,-12,-19,-15,13,16,10,9,14,7,15,-4,9,7,-8,-13,-9,1,11,-2,-21,0,13,-6,6,19,16,0,-2,0,1,11,15,0,-8,8,-1,-9,3,15,22,-4,-15,-11,-13,-11,-15,0,-4,14,5,-1,-4,7,3,-11,-3,3,-5,-13,-22,4,1,16,9,7,0,0,0,-7,-4,-6,-6,-15,-3,-4,-12,0,-1,-10,-6,-9,-21,-16,-4};
 
localparam signed [width-1:0] weight [0:output_number-1][0:input_number-1]='{
{-6,-14,-1,1,-1,-12,-7,-67,-4,-9,2,3,-21,-5,-523,-37,4,-8,-4,-1,-7,-2,6,-33,-19,-106,-16,5,-1,-11,-8,-23,-7,-6,-26,-82,-64,-187,0,0,-13,-5,-2,-36,-7,-11,-14,5,-5,-11,-4,-6,-88,-10,-8,-17,-5,0,-5,-1,-12,-4,-1,-58,-53,-37,-4,-14,-11,-5,-6,-11,-15,-6,-12,-1,-15,-9,-16,-19,8,-72,-3,-34,-63,-14,-1,-8,-14,-5,-39,-2,-23,-8,-15,0,-11,-5,-12,-17,-6,-26,-17,-12,0,3,-9,-16,-289,0,-1,6,-17,-16,-8,-103,-6,-7,-11,-44,-9,-5,-3,-9,0,0,-20,-7,1,-2,-7,-58,-3,-1,-11,-1,-14,6,3,-2,4,2,-12,-15,-7,-10,-10,-6,-23,-11,-3,-4,0,-142,-2,2,-11,-10,-7,-11,-3,-7,-13,3,-77,-3,-14,-3,-12,2,-29,-9,-15,6,-3,-9,-14,-3,-8,-7,-14,-34,4,-14,-111,-4,1,-9,-17,-22,-2,-36,-26,-10,-1,-18,-16,-24,-3,-3},
{-2,-1,-3,-8,-3,-6,6,-58,-16,-11,7,-8,-25,1,-517,-34,7,-16,-9,5,6,-5,0,-18,-12,-125,-4,-2,-10,-2,0,-20,0,0,-24,-81,-70,-199,-4,2,-7,0,-15,-44,-8,-13,-7,-9,-4,-5,-19,-11,-66,-14,-2,-10,-5,0,-12,-1,0,0,-8,-47,-63,-45,-6,0,-3,-14,-19,-17,-5,5,-2,-10,-13,-17,-9,-17,7,-65,0,-26,-52,1,-1,7,-1,-4,-35,0,-27,-8,-9,0,-12,-18,-10,-1,-7,-18,-13,-15,-2,4,-6,-11,-240,1,-11,1,-1,-18,-1,-116,-10,-15,-4,-42,1,-11,2,5,-14,-1,-18,0,-6,-2,8,-70,5,-2,-10,-7,-3,-4,6,6,-3,-8,-2,-14,-15,-1,-12,0,-31,-13,0,-10,-7,-173,-14,5,-2,-12,-16,-18,-9,1,-8,-3,-82,6,1,1,0,-7,-26,-15,-9,-6,7,-13,-11,-12,-7,-10,-14,-40,0,-4,-125,-14,-14,-19,-14,-9,-3,-36,-17,-14,-3,-14,-14,-18,-7,4},
{-4,-526,8,-25,5,-10,-3,-2,-21,-11,-5,20,-109,-47,-96,-25,-21,-38,-4,1,-3,3,6,-15,-129,-12,-17,-5,-129,-16,4,-12,-5,-28,-15,-20,-12,-70,-21,-3,-3,5,9,-26,-23,0,-77,6,5,-15,-10,14,-2,-16,-26,-364,-42,-2,2,-7,-11,14,-25,-29,-537,-23,-6,10,0,-11,-8,-10,-11,8,-11,-7,-19,-10,-10,-424,3,-180,-9,-9,-72,12,-46,0,1,-14,-44,1,-6,-10,-6,-260,-18,-5,18,-14,-884,5,-20,4,6,-5,3,16,-47,-6,7,0,-11,-17,-11,-81,-3,0,-30,-29,-16,-34,-106,8,-7,2,-7,4,-12,4,7,-17,-3,-33,-20,-2,-129,3,-8,6,8,-128,-9,0,-5,-12,-13,-7,-14,-3,-81,-8,2,-33,-16,-6,17,-8,-3,-19,3,0,12,7,-27,0,14,-32,-25,0,-10,-6,-84,-9,-8,-15,-3,8,-1,5,-13,-15,-6,-1,-30,-14,-37,0,-22,-44,-313,-19,-13,2,-6,-171,-10,-16,-1,-29},
{-11,-75,1,1,13,-14,-6,17,0,-161,2,50,-154,-3,-64,-75,-3,-4,0,-8,-10,2,-6,6,0,-2,-37,-9,11,-38,-1,22,4,-53,0,9,-12,-33,3,-56,-65,4,9,-38,-26,12,0,-7,-2,16,10,14,-62,1,-25,-102,-1,-7,-6,-13,-51,-257,0,-4,-75,-20,17,8,23,-105,-8,-36,2,-8,-609,-26,-14,4,-2,-514,-1,-40,-57,-86,-9,7,-45,-2,-2,-258,-99,-4,-1,0,-107,-303,-17,22,34,-56,-80,-4,-60,14,3,3,6,15,-3,9,13,-25,-21,39,-3,-71,-4,-44,-48,-20,-60,-19,-92,27,-10,3,14,-13,6,0,-2,-1,4,-6,-32,-35,-24,3,-6,6,-1,-47,5,-39,21,-74,12,-19,-93,-55,-92,19,-3,-16,10,-3,27,-613,-12,-18,-4,8,19,0,-41,-2,21,19,-95,15,15,-6,-136,4,0,7,-17,-5,-3,10,8,-30,-6,-188,-18,-56,4,-475,-205,-188,17,6,-14,19,2,13,-17,-39,6,-915},
{-19,-47,0,-12,2,-1,6,6,-1,-116,-2,24,-59,-8,-74,-20,6,-13,0,-6,-3,0,-9,4,0,4,-41,-3,16,14,2,16,29,-34,-7,4,4,-19,7,-38,-20,-2,25,-49,-42,16,0,-6,-1,12,-11,15,-9,11,-10,-14,-6,-2,0,-18,-12,24,1,-5,-236,-12,10,-12,11,-447,-17,-64,-10,4,-26,-28,-5,4,-9,-545,0,-88,-49,-18,-20,17,-26,3,20,-525,-21,-6,-12,-7,-108,-129,-11,7,6,-51,-900,-10,-27,17,7,4,13,6,-5,5,13,-23,-24,18,3,-57,-14,-25,-55,-16,-46,-16,-9,39,-6,-5,1,-20,13,-2,4,5,4,2,-58,-18,-9,2,-1,0,-1,0,-1,-41,13,-43,15,-7,-130,-40,-34,14,3,0,3,-6,26,-43,-10,-17,-5,2,5,-8,-25,-8,21,12,-78,33,21,0,-20,1,2,-2,-4,-4,5,26,32,-74,5,-13,-9,-37,-372,14,-323,-128,-519,5,1,14,7,-116,0,-9,0,-33},
{-15,-46,0,4,0,9,5,0,0,-49,8,46,-144,-31,-59,-22,-7,-12,20,-7,4,2,-1,-5,-29,3,-112,2,-37,-11,-4,22,-34,-14,-27,17,4,-16,0,0,-6,3,10,-26,-18,14,1,0,-4,-18,6,13,22,0,-40,-63,-14,-3,-9,-7,-8,59,0,-7,-285,-14,-3,-8,-4,-384,-12,-55,3,-4,35,4,0,-6,-3,-617,-2,-35,-10,-3,-27,20,6,2,-24,-597,-33,-13,-10,-5,-17,-125,-19,26,37,-47,-111,-27,-20,4,-2,-6,-12,27,-2,-6,15,-25,-32,18,-9,-33,-6,0,-37,-31,-24,-9,-46,26,-16,3,-13,-2,-6,4,8,-4,-7,-2,-53,7,-59,-2,3,-9,-2,-25,4,3,19,-12,-18,-3,-150,-16,0,22,4,8,2,-1,17,-291,-6,-17,29,5,-4,-1,-34,-8,10,-27,-22,20,18,-3,-45,1,6,-36,-11,14,-8,-8,-7,-51,-5,-17,-2,-14,-177,53,-139,-109,-158,17,-9,8,5,-205,-9,-17,0,-52},
{-29,-65,-4,4,2,5,-4,4,-14,-28,-6,22,-146,-45,-37,-20,12,-14,26,5,-5,-10,3,-27,-18,-5,-251,1,-73,-26,4,-6,-48,2,-36,7,-8,-23,2,5,-8,3,12,-39,-13,10,-11,-2,7,-24,-7,26,19,-17,-51,-45,-3,-5,-19,1,-13,60,13,-15,-187,-18,-8,3,0,-319,-9,-27,0,0,43,14,-16,-23,-10,-580,-2,-2,7,8,-32,3,0,-8,-16,-773,-46,-12,-13,-11,-12,-176,-16,12,27,-27,-145,-11,-8,3,-8,-3,-19,24,-11,-8,15,-7,-34,5,-7,-56,-9,8,-38,-29,-8,-5,-32,20,-1,-6,-14,7,-18,0,0,-2,-1,-26,-26,-3,-81,-6,-1,-8,3,-65,-12,19,2,11,-36,-8,-95,12,10,9,0,0,13,-6,24,-759,-11,-24,34,3,-1,-6,-39,8,13,-106,-16,11,0,-22,-51,0,0,-31,-8,32,0,-11,-23,-2,-2,-58,3,1,55,41,-84,-100,32,3,-7,-1,0,-157,-3,-6,7,-32},
{-92,-27,-1,-7,-1,4,-10,9,-26,-19,5,34,-97,-39,-22,-457,2,-19,37,-4,-1,-2,-7,-18,-32,-10,-63,-2,-89,-31,1,-13,0,-11,-27,10,4,-26,-20,0,-21,-1,27,-1,-18,5,-9,-2,2,-21,-27,14,8,-15,-4,-21,4,3,-6,40,-19,35,56,-10,-88,-20,-20,4,-6,-13,-33,-27,-19,-3,14,0,-12,-40,-8,-850,-5,-9,3,-5,-38,14,-7,6,-14,-637,-63,-3,-13,-4,-7,-711,-15,14,9,-5,-45,-20,-6,2,4,0,4,23,-13,-23,1,2,-12,-22,-7,-147,-54,17,11,-18,-15,4,-5,22,-1,-3,-5,18,-15,-8,-10,-4,0,-38,-13,-8,-29,5,-8,5,-7,-59,-7,12,15,3,-23,-9,-52,10,-14,-3,2,-8,2,-13,16,-35,-6,-24,35,7,-17,3,-23,-3,13,-4,-8,16,-4,-15,-29,-1,3,-20,-23,36,0,5,-9,-5,-9,-116,-5,-19,-7,13,-25,-53,-15,16,-19,-11,-9,-53,7,-11,6,68},
{-166,26,-5,-17,5,5,-6,23,-24,-9,-10,22,-89,22,-21,-235,-8,7,-22,3,4,-9,5,-25,-55,-3,-17,0,-66,-6,-3,-21,-12,-27,-22,-4,14,-14,-33,-2,-8,-4,11,-47,-29,4,1,5,3,-12,-9,-4,-3,-16,-13,3,2,-4,-18,45,-19,-10,47,-3,-57,-1,-19,12,-6,-3,-86,-7,-32,2,-50,0,-12,-87,-18,-614,8,-33,17,-17,-114,-1,-15,7,-9,-261,-85,0,-18,-8,-19,-412,-9,11,23,4,-52,-9,-17,-14,4,-8,0,-16,-66,-2,0,-1,-7,-13,0,-171,-202,14,3,-26,0,-18,5,22,-67,-9,3,10,-18,-8,-3,-4,-10,-105,-15,-13,-13,-5,3,6,-1,-37,-2,18,13,15,-18,-21,-38,-26,-105,0,-2,-7,-4,-13,-8,-18,-10,-21,-77,0,-11,6,-3,0,7,84,-18,21,-3,-16,-72,-1,-7,-2,-76,-8,-4,7,-19,-4,-4,-147,-17,-11,-9,13,-24,-55,-26,1,-14,-24,-3,-16,25,-17,-2,-33},
{-251,6,-8,-12,-5,-8,-8,12,-13,-1,-4,14,-116,0,-3,-318,-9,4,-19,6,-5,3,-7,-20,-80,-13,-20,4,-44,2,2,-14,1,-18,-6,-11,7,-16,8,-7,9,0,-35,-44,-7,8,7,-7,-2,-3,0,-20,-19,2,-19,-48,-2,2,-1,-190,-9,-70,-26,-7,-40,-35,-4,-10,-1,6,-113,1,1,7,-31,-2,-16,-109,-4,-73,8,-51,-4,-27,-219,7,-10,-3,-2,-639,-87,-8,-16,-2,-3,-17,-6,-10,21,4,-7,-78,-54,1,-1,-2,-2,15,-127,-6,-10,-7,-9,-3,-10,-62,-17,-6,-5,-22,10,-2,-39,14,-12,0,-8,0,0,-5,-10,-22,1,-118,-1,-11,-38,0,-9,7,6,3,-4,8,3,0,-9,-18,-33,-31,-57,0,6,0,-6,-7,-36,-18,4,-8,-69,2,2,2,-16,-7,-3,41,-12,6,10,-6,-39,2,0,-4,-17,-54,-7,-9,-13,-3,3,-331,0,-5,4,3,-26,-48,-6,5,-25,-41,5,-9,-113,-5,2,-37},
{-252,-4,0,0,-25,-15,-2,10,-1,5,-1,19,-89,4,-7,-373,-20,-9,-11,-3,-7,-8,-2,-5,-51,-3,-6,0,-4,0,-1,-20,-1,-12,-15,1,-2,-23,-3,-15,-5,-2,15,-33,-6,0,5,3,-2,1,-14,7,-66,1,-8,-169,-23,-7,-6,-16,-21,-7,-15,-4,-55,-55,-17,19,-1,4,-59,-12,3,-8,-19,-11,-9,-64,-6,-74,-4,-61,-6,-53,-371,4,-7,0,7,-328,-73,-7,-10,-1,-4,-209,-10,-5,8,-18,10,-25,-23,-7,-8,-9,-2,-23,-170,-8,5,5,4,-15,2,-147,-10,-5,-12,-29,-2,-9,-118,15,-27,3,0,-26,-7,1,-9,-170,-5,-25,0,-4,-20,-1,7,5,6,-3,2,-22,1,0,3,-8,-24,-10,-37,-6,1,-21,-10,-11,3,-96,-20,-11,-21,-8,-7,-5,-21,-5,-16,7,-7,6,11,-6,-33,-1,3,-6,-13,19,4,6,-1,1,-3,-263,-5,-17,-20,-44,-18,-35,-38,0,-17,1,-1,-3,-72,-53,-3,5},
{-41,-12,2,16,-9,-12,-5,1,-13,3,4,21,-53,-14,-17,-247,-20,-5,24,-7,3,1,-8,-3,-73,7,-9,-4,-28,-3,3,-7,-3,-2,-28,-2,-3,-25,-5,-8,10,-5,5,-42,6,-14,-8,-6,-5,-12,-24,-34,-48,-2,-18,-38,-2,-4,-8,-37,-37,5,-12,-32,-49,-40,-31,-8,10,0,-10,-24,3,3,-18,6,-3,-28,-6,-497,0,-122,1,-38,-102,-12,2,2,-3,-66,-45,0,-9,-7,3,-347,-15,-5,4,-53,10,-38,-10,-41,0,-8,1,18,-45,-19,-2,-19,11,0,-8,-135,-8,-18,-2,-28,-19,3,-360,10,-2,5,-2,-9,-9,1,-4,-14,-3,3,-19,-31,-17,-5,0,-4,-3,-27,-4,7,-5,1,0,-14,-23,-11,-14,-26,0,-20,-9,-2,5,-82,-22,-41,15,-2,-5,4,-36,2,-50,-115,10,-12,5,-1,-37,5,-1,-5,-16,22,-2,-4,-7,-20,6,-420,-10,-26,-41,-42,-8,-9,-54,-13,-27,-9,-1,11,-61,-23,2,19},
{-14,-14,-1,-2,-3,-3,5,-62,-9,-3,4,-1,-16,-6,-503,-35,-2,-4,-11,-3,-4,6,3,-35,-6,-125,-12,-4,-5,0,-3,-14,-1,-3,-18,-79,-60,-162,-11,-14,-10,-5,-3,-46,-11,-10,-13,-3,2,-1,-17,-13,-72,-12,0,-15,-10,-2,-4,-10,-3,1,-4,-50,-57,-47,-7,-17,-4,-11,-6,-16,-4,3,-11,1,-29,-6,-5,-16,-7,-78,0,-31,-50,1,-1,-7,-14,-15,-40,-12,-30,6,-12,-14,-20,-12,-14,-3,-1,-26,-28,0,-9,6,1,1,-212,-11,3,-4,-1,-6,0,-117,-4,-6,-12,-34,-14,-10,-14,4,-5,-1,-13,-3,0,-7,-3,-68,5,-17,-4,-1,0,-5,-7,1,8,0,-5,-16,0,-14,0,3,-29,-9,-7,-1,2,-184,-5,-1,-13,-8,-3,-29,-14,8,-8,6,-83,7,1,-1,-4,-13,-20,-17,-13,-4,2,-7,-8,-15,0,-17,-6,-42,-3,-10,-130,-8,-9,-20,-21,-21,-13,-45,-15,0,3,-8,-20,-23,4,-6},
{-2,-14,-1,-14,0,-1,-1,-63,-10,-13,-2,1,-18,-8,-516,-41,0,-13,-12,-5,-7,6,-7,-31,-6,-113,-13,7,-4,-9,6,-10,-6,0,-14,-72,-66,-179,-2,-13,0,-8,-14,-48,-5,-7,-13,3,-4,0,-12,-11,-77,-5,-1,-17,-14,5,-1,-8,-13,-13,-12,-51,-59,-53,-10,-10,-1,-1,-14,-10,-10,5,-12,-4,-30,-7,-13,0,8,-79,-6,-29,-55,-10,-15,4,-13,-4,-30,-2,-18,0,-1,-1,-20,-16,-3,-11,0,-27,-15,-4,7,-3,-14,-6,-263,-2,-11,0,-9,-10,-10,-115,-11,-11,-10,-47,-14,-1,-3,-5,-2,7,-7,-12,2,-2,0,-65,-2,-1,-15,-3,0,0,6,3,-5,-8,0,-11,-13,-7,0,-4,-26,-19,-17,-6,-9,-170,-12,-1,1,-19,-14,-22,-11,4,-1,-2,-90,0,-8,1,1,-14,-43,-20,1,5,4,-4,-6,-5,-10,-13,-5,-32,0,1,-111,1,-2,-20,-9,-15,-10,-30,-12,-13,5,-11,-3,-20,0,5},
{-1,-4,-5,-7,-10,-3,-4,-77,-10,2,-6,0,-27,-11,-510,-44,-7,-12,-1,0,3,-7,-8,-41,-10,-111,-4,5,-15,-14,-4,-15,-1,-17,-19,-69,-63,-169,-4,-15,1,-5,-8,-45,-8,-11,-7,-1,1,-11,-8,-9,-82,-10,-16,-17,-12,-7,-16,-8,-14,2,-14,-52,-53,-35,-8,-1,-2,-13,-6,-10,0,4,-9,0,-26,-11,-12,-13,-7,-69,-11,-28,-51,-12,-1,1,0,-6,-28,-16,-16,-6,0,-5,-18,-2,-10,-8,-4,-31,-26,-10,5,1,-12,-15,-281,-12,-13,-2,-6,-12,2,-96,-2,-1,-20,-36,-5,-12,2,-2,-3,2,-16,-5,1,4,0,-61,3,-15,-9,-8,-13,-4,6,-7,0,-13,1,-2,-4,-12,-4,0,-25,-17,0,-4,0,-169,-13,-4,-6,-7,-1,-21,-4,1,-5,4,-82,-7,-1,-2,-5,-12,-38,-11,-7,0,5,-2,-13,-10,-9,-9,-11,-42,4,1,-118,0,0,-10,-11,-13,-3,-34,-20,-2,-5,-19,-14,-20,-3,-8},
{-62,0,-6,-11,11,19,0,9,-8,-18,-5,0,-16,11,-31,-161,-15,-10,-44,2,3,7,6,-31,-39,-10,2,5,-10,4,1,6,-4,-5,-21,-12,-13,-50,-1,21,15,-2,-7,-22,-10,4,-13,-1,-6,-13,-18,5,-27,-16,3,-31,-18,0,-9,11,1,-34,8,-36,-37,-9,-10,25,0,0,-409,-28,0,-3,-22,-11,-10,-56,-29,-51,1,-42,13,-12,-34,7,-38,-7,6,-69,-49,-2,-8,4,-23,49,0,0,18,-3,-6,-111,-26,14,-6,-5,-13,-23,-229,2,-21,0,-17,-2,4,-249,-21,16,5,-30,4,14,5,5,19,2,-30,7,-16,-1,-4,-31,-3,-292,-15,7,0,6,-5,2,0,5,-9,10,-9,-3,-25,-18,0,-50,-13,-11,-7,-35,-9,-8,-80,1,2,-4,-100,3,6,3,-40,6,11,15,-15,17,-3,-11,13,5,6,-5,-29,-52,4,-25,2,-21,2,1,-27,1,-2,3,-8,7,-4,-1,-16,-25,0,-33,-231,-91,0,-8},
{18,-25,6,-28,-18,-13,-10,5,-3,-31,0,-22,-40,-7,-40,-659,-17,-27,-34,5,6,-7,-8,-15,-7,8,-17,-3,1,4,-2,-16,-22,-11,4,8,-18,-25,-13,-21,3,0,-5,-46,-17,23,0,-6,-2,-18,-8,-4,-5,-18,16,-2,-27,5,-12,-7,-61,-4,-14,-48,-82,-11,0,-12,-3,-18,-21,7,-35,0,-4,-12,-307,-52,-3,-128,6,-35,0,-4,-6,-2,-19,8,18,4,-31,-1,-11,4,-39,-6,-11,-35,2,0,10,-59,-35,-18,-5,-2,1,-6,-15,-27,-18,0,-10,-8,-3,-837,0,-38,17,-23,-6,0,5,-3,-143,2,0,-1,-5,-4,-1,-3,-3,-16,0,4,6,2,-8,-9,-3,-20,-1,-3,-16,0,-28,-10,-24,-21,-16,0,-6,-8,-18,-6,0,-138,-6,-18,-5,0,21,2,-10,7,-1,2,-12,-27,0,-1,-19,-7,-7,-21,-419,-20,-4,10,10,8,-5,-91,0,6,-3,-88,-21,-29,-40,-16,1,0,-9,-9,16,-4,-10,6},
{30,-53,5,-34,4,-24,-6,8,25,-86,-6,-99,-38,-17,-49,12,-9,-34,-42,8,-7,4,0,0,19,16,0,-11,0,7,1,-11,32,-26,25,34,-19,-3,-7,-34,-5,8,7,-23,-46,12,-22,-1,-10,2,-13,8,-3,16,37,15,-20,-1,8,0,-47,-30,6,-23,-107,-16,38,-5,-10,-125,-9,-4,-20,-11,15,-29,42,27,24,-251,6,-49,-10,-32,-8,7,-47,-2,31,-14,-14,-103,3,-10,-98,-67,-6,-64,-27,-37,25,-35,-57,2,-2,-3,-30,-10,-29,2,-36,7,-11,4,-11,2,10,-17,13,-10,-17,-13,9,-31,-3,-2,4,-16,21,-9,-4,3,0,-1,-1,-7,-1,-2,-5,6,7,-34,27,-25,-23,-22,10,-19,-39,-29,-52,0,1,7,-19,-4,20,-92,-2,-10,-34,-3,7,-5,21,1,29,6,-25,21,13,1,32,0,-2,-5,-15,-24,-8,5,37,19,4,-65,14,-12,-31,-32,-129,-36,-36,-37,7,27,-3,-23,4,-24,-3,19},
{5,-28,-8,-43,24,-16,-2,22,11,-35,-2,-150,4,-13,-49,-11,2,-35,-19,8,6,0,-14,18,14,9,-12,-4,10,24,0,8,29,-46,0,49,34,1,-10,-29,-18,6,4,-12,-38,3,-13,7,-6,7,-1,-4,22,14,21,8,-34,-8,0,-36,-29,-64,-32,8,-82,-9,16,-6,-16,-20,-23,-23,-36,-3,36,-27,25,34,7,-128,8,-26,-22,-4,-8,-18,-29,-2,8,-32,2,-103,8,6,-71,-156,-10,-78,12,-56,34,-6,-47,-19,-4,3,-29,11,-30,8,-36,-8,-11,5,-10,13,-23,-24,8,-7,-30,-33,13,-60,-106,-3,-10,-11,18,4,-3,18,-8,36,-20,-14,0,-1,-1,1,-5,0,6,-27,-22,-36,39,-19,-92,-13,-38,12,-7,11,-8,-13,10,-135,-4,-18,-17,5,3,1,6,-3,104,6,-23,11,22,6,-38,-4,-1,19,0,-4,7,-16,46,6,0,-95,26,-20,-11,-85,-126,-34,48,-17,10,15,0,-19,-15,-12,0,31},
{-81,-53,4,-7,12,3,-3,33,-16,-24,3,-129,-39,-39,-28,12,-1,-24,42,-4,5,4,-3,0,1,11,-216,-2,-45,11,6,11,-58,-18,-35,30,25,-1,-17,8,-32,5,39,-27,-15,20,-11,0,-5,-35,18,13,52,-12,-31,-14,-17,0,-32,-19,-14,87,-15,5,-118,0,-1,4,-14,-43,-46,-40,-7,-7,30,8,30,6,28,-24,0,6,-21,12,-1,9,-18,-8,-4,-41,-28,-171,21,6,9,-74,-10,-65,16,-28,27,2,-23,0,-2,-8,-35,46,-23,-4,-21,-1,-17,-5,-9,13,-29,33,-15,0,-5,-11,15,-39,-9,6,-9,10,-27,-6,-9,15,3,26,-67,12,-40,4,3,-9,1,-17,-4,4,-6,-7,-18,-10,-114,27,12,7,-2,9,16,-10,16,-19,4,0,35,-7,15,-5,-16,0,64,-14,-51,6,17,6,-98,5,-3,-41,46,22,-1,-15,39,17,-10,-39,16,-6,-26,-8,-138,-16,52,0,-4,-1,-14,-173,10,4,-3,37},
{-188,-41,4,17,6,16,1,32,-51,-17,7,-123,-40,-61,-20,27,1,-1,57,-8,-5,3,-10,-23,-9,-1,-193,-8,-73,-19,-1,-13,6,-10,-36,25,18,-6,-6,16,-4,0,30,-58,-4,30,-18,-6,2,-43,-3,23,53,-21,28,-15,0,3,1,24,4,48,22,16,-117,1,-30,2,-13,-79,-59,-21,2,-11,-26,5,28,0,20,9,-5,8,0,5,7,30,-20,-1,-11,-62,-18,-57,14,-5,31,14,-8,-57,20,-7,-76,14,-15,-8,1,6,-22,42,-25,-23,2,1,-28,-15,3,-4,13,29,26,-6,2,7,1,-21,-10,-1,-5,25,-44,2,-11,-7,-5,-10,-42,15,-36,3,4,-4,1,12,-4,29,1,0,-33,7,-63,29,13,15,-4,13,3,-3,7,-93,-7,-12,48,0,1,1,-35,-4,61,-18,-32,-19,11,1,5,-8,4,-34,11,45,-10,-14,38,30,-5,-15,19,-5,-52,-4,-82,-39,60,20,2,-27,-8,-149,-41,-13,-7,20},
{-235,51,6,16,-6,21,-1,44,-45,-19,1,-51,-20,-7,-11,21,-1,12,10,0,-5,0,-4,-10,-16,-1,31,-1,-84,-48,1,-10,20,-7,-18,18,21,-12,16,22,-11,-6,7,-66,23,11,-21,-6,0,-16,-2,19,43,-15,39,-10,17,3,40,65,63,-73,86,23,-64,-14,-24,39,-28,-44,-77,-4,-1,-3,-99,-2,13,-15,23,14,-1,11,28,2,-19,9,-23,-3,-18,-74,-38,-166,16,-9,43,17,-10,-15,28,-13,-215,-11,-47,-35,3,-1,-16,-38,-4,-14,20,-4,-18,-22,-5,-4,16,4,19,-21,2,-10,1,-13,-21,-2,-10,8,-15,3,-8,-35,-2,-9,-16,-17,-2,5,5,6,0,95,-2,14,27,11,-9,-3,-32,-12,6,10,0,1,-1,-6,-2,-117,-15,-8,-39,5,-21,-5,-18,8,45,34,0,9,11,3,-34,-4,-3,-3,-6,33,-4,-15,17,31,2,-115,13,-13,-47,-82,-16,-39,25,25,-2,-17,2,-15,-44,-82,1,0},
{-179,102,-1,30,8,45,8,24,-35,-16,-9,27,-18,43,22,-16,-7,13,-47,3,-3,5,0,0,-23,-18,5,-5,-31,-11,-6,6,-12,-10,-6,16,21,7,18,36,2,5,-60,-118,9,1,-18,6,5,-18,-3,9,26,-36,-16,0,15,0,14,46,52,-5,60,24,-32,-15,-22,12,-46,8,-80,-12,5,-8,-53,-45,21,23,23,20,-8,-7,56,-15,-34,4,24,-8,-19,-67,-52,-31,3,3,26,64,-9,11,30,0,-74,-4,-72,-44,-7,8,-24,-60,28,0,25,1,-7,-8,-9,-1,-25,-40,-106,-11,2,-21,18,-1,0,3,6,-14,-7,1,-7,-39,3,-17,5,-13,-15,8,-4,3,-3,72,1,-4,39,3,-6,-1,-19,-78,-31,13,-6,18,18,-5,-51,-54,-21,-4,-122,8,-30,1,4,4,-3,44,5,-9,15,1,-54,1,5,-11,9,-71,-7,0,-8,35,-1,-141,21,-5,-14,4,-32,-41,-7,32,-11,-31,-12,15,-60,-97,-5,-111},
{-131,77,-5,19,-35,20,0,32,-19,11,-12,26,-7,20,15,-51,-15,20,22,8,4,5,-11,-6,-36,-9,-37,0,24,0,3,-31,-17,-5,-6,12,21,4,-14,1,28,8,-67,-78,1,6,-21,-2,-3,-2,12,-10,-13,-15,-18,2,18,5,-15,-42,-4,44,-68,14,-3,-60,3,-48,-26,0,-33,6,-4,-5,48,-57,0,6,33,20,-5,-3,1,-16,-26,12,27,-3,-10,-43,-41,35,43,4,1,79,-11,28,35,-30,-20,15,-34,-12,-7,1,-28,-3,29,8,12,-12,-24,18,4,29,-61,-24,-111,2,0,-1,4,19,12,-5,0,-75,-13,5,-3,-7,-6,-52,0,-18,-17,1,-5,1,0,6,-10,-69,28,-50,-7,1,-16,-57,-23,21,-7,7,-13,-7,-33,14,-33,-2,-7,6,-40,-4,3,-6,-78,-33,-1,-66,11,1,-47,2,0,13,39,-42,-4,-9,-19,36,-5,-161,20,17,26,38,-51,-28,-18,33,-10,-25,-3,-3,-120,-36,4,-45},
{-97,28,5,4,-63,-35,5,32,-11,9,4,26,-4,-14,5,-86,-4,14,-1,4,-9,3,-12,-4,-42,-10,-45,-10,2,33,1,-52,-4,-15,-5,-4,12,-4,-11,-34,13,-3,20,-63,-4,-10,-6,5,3,-2,-29,-46,-25,0,-16,-15,28,4,-8,-100,-46,17,-64,12,5,-45,13,-3,-4,-7,-11,2,-29,0,77,-35,-24,7,30,0,-6,6,-5,-5,-22,-15,-3,-6,7,-36,-46,58,75,-5,-2,83,-10,23,40,-66,-5,-1,-2,-56,-6,-7,-17,-10,10,17,4,6,-20,10,2,16,-98,32,-44,-4,-24,-5,0,22,16,3,12,-34,-17,-5,0,14,6,-87,-1,-50,-20,3,4,-4,-1,-22,-15,-40,23,-18,4,6,-5,-52,-13,22,4,8,-47,-19,17,15,-112,-14,23,0,-14,0,5,2,-130,-82,8,-34,-11,-1,-41,-8,-3,0,46,41,6,-5,-21,23,2,-95,21,-28,19,21,-29,-21,-23,21,-23,-1,0,-3,-123,-17,-7,0},
{-107,-14,1,-21,-30,-27,4,26,-27,-1,-7,35,-9,-32,28,-143,-6,-17,12,0,2,-5,-10,-2,-27,-6,-18,4,-28,21,-7,-8,5,-23,-2,-8,8,-2,0,-29,-2,-6,29,-57,21,-11,-29,-10,4,-5,-102,-42,-43,0,-22,-9,8,7,-11,-108,-51,-37,-50,6,-5,-46,0,6,7,-15,-15,4,-14,-10,35,-17,-79,2,40,-14,-4,-24,11,28,2,-14,-8,-2,11,-22,-35,61,79,-1,-2,18,-23,4,25,-64,11,-1,-17,-125,-2,-4,-17,34,-5,0,-9,-3,-19,6,-5,29,-123,78,-28,-36,-24,-11,-4,20,13,-3,13,-20,-6,1,-7,18,6,-138,8,-67,6,-3,0,5,2,-50,-19,-2,7,-15,-7,-1,8,-34,-28,22,-7,-13,-49,-19,27,17,-93,-39,18,-4,-7,-8,3,-6,-77,-66,8,14,1,-26,-14,-3,3,-10,61,30,-9,0,-19,17,-8,-14,5,-92,-16,40,-18,-1,-36,12,-21,18,0,-13,-88,-15,-8,20},
{-103,-20,8,-26,-13,-45,-8,18,-20,-13,-6,30,-1,-41,21,-129,-8,-13,7,-2,-2,-1,-13,1,-9,-14,-28,0,-29,22,-6,11,0,-1,-20,0,5,-6,-4,-38,1,3,31,-53,2,-21,-38,2,4,1,-117,-24,-52,2,-14,3,13,-1,-24,-102,-36,-38,-36,-6,-8,-40,2,-49,7,-10,-16,-4,-5,-10,-18,35,-105,21,13,-28,-7,-45,-13,-5,0,-20,17,2,-8,-66,-14,57,56,-9,-6,-74,-7,5,23,-89,11,-10,-54,-185,7,-7,-23,13,-53,-3,-6,-11,-28,8,-8,47,-124,44,-17,-27,-43,-13,-6,20,18,4,-8,-11,-3,-2,3,40,-3,-86,7,-60,10,3,-10,-9,-2,-61,-21,18,11,13,-5,-3,-5,-34,6,16,-6,-30,-24,-8,20,12,-63,-37,15,2,-15,4,-6,4,-117,-12,11,7,-3,-35,3,1,2,-5,31,1,-4,-8,-1,6,-3,15,-23,-110,-21,46,-26,-2,-13,11,-20,14,2,-6,-46,10,2,0},
{-38,-17,-7,-31,-22,-11,-5,-3,-2,10,-5,20,-19,-86,-19,-12,5,-672,-14,8,0,3,0,-5,5,-85,-21,-3,-34,2,6,-51,-1,-6,-7,-44,-10,-41,-18,-4,7,4,-15,-92,-5,5,-6,-2,-5,-3,-21,12,-619,8,-54,-6,7,-9,-14,-328,13,0,-132,-16,-24,-766,10,-96,1,-19,-19,-16,-9,-4,-2,-10,-59,7,5,-33,5,27,-31,-43,-29,4,-29,-3,1,-18,-2,-4,-2,-4,20,-14,-10,0,16,-20,9,-290,-152,25,1,-7,-7,-1,-73,-14,-3,-12,-6,2,-2,-103,-21,-12,-68,-60,-67,-97,1,9,-29,3,-2,-27,3,0,0,-55,-6,-234,10,9,-10,8,-6,3,-3,-210,27,-23,-4,1,4,-24,-60,-22,-36,-1,-9,-31,-24,4,-21,-10,-59,3,-1,4,-4,3,-9,-3,-2,-19,8,-136,-28,13,-18,3,-2,-11,0,-175,4,1,2,4,-7,-10,-12,32,-6,-59,-12,-631,-13,-6,-22,1,-5,0,-22,-43,7,4},
{-17,7,-1,-6,-278,-14,0,0,-5,-2,0,-17,-28,1,-90,-269,-9,-4,1,-6,7,6,-7,-24,-4,-967,-14,-6,3,-48,0,-17,-339,-18,-10,-7,-6,-57,-150,-12,-8,0,-1,-55,-9,3,-53,5,0,-7,-9,0,-1,-122,-24,-12,-8,-5,-40,-8,-5,9,-431,-15,-25,-31,0,-11,-7,-229,-100,-3,-33,8,2,-9,-10,-157,-14,-357,0,-4,-10,-65,-42,6,-19,0,-10,-4,-26,-6,-23,-10,-8,-5,-13,6,21,1,-371,-20,-28,-275,4,-3,-10,-21,-154,-8,-10,-7,-68,-8,5,-262,-281,-33,-150,-37,-5,-14,0,12,-5,-7,-14,6,-19,4,1,-417,-5,-11,-4,7,-4,7,-7,-1,0,7,-29,-12,5,-8,-54,-16,-70,1,-16,9,-1,-33,0,1,-7,-14,-110,-15,-3,3,-4,0,-8,4,7,0,-15,-20,12,-343,-14,7,1,-293,-257,-8,4,-19,-9,4,0,7,-41,-11,-12,-4,-12,-34,9,11,-13,-18,-6,-8,-7,-97,0,-11},
{33,-13,7,-22,-40,-12,-20,-10,20,-10,-9,14,-10,8,-32,0,-17,-19,-37,3,-4,2,-5,-23,21,0,-79,0,13,-22,0,-31,-19,-5,13,-6,-7,-39,-21,-27,2,-3,9,-41,-22,9,-24,-10,5,1,-7,9,-93,-2,-8,4,-19,-9,-30,-34,-10,-71,-101,-14,-58,-9,14,-2,7,-65,0,0,-28,-6,-6,18,22,-15,18,-66,0,19,-8,-19,-21,14,-5,-8,4,25,-27,-671,28,5,3,34,-29,-13,18,15,30,-33,-43,4,4,1,-28,-11,-49,-33,-24,-22,-2,-14,-2,-17,-28,-20,-51,-26,-45,1,5,3,-45,0,-17,-5,0,0,-7,-9,-1,-56,3,25,-2,-2,-1,6,-5,11,-12,-6,-25,-26,-6,-16,17,16,-16,-13,4,-15,-24,-19,-9,-44,2,10,-28,3,17,5,-4,-6,-116,0,11,-11,-2,-8,-19,0,3,5,-1,-15,0,1,14,-21,2,-39,17,10,32,-27,-36,7,-64,-18,-1,-15,3,-12,-8,44,-9,-3},
{23,-24,-4,-32,-56,-12,-5,-40,24,-19,-4,9,-7,2,-57,24,-20,-25,-56,-6,-4,3,-3,11,6,2,-21,0,15,-16,-4,-5,-1,5,28,27,-7,-4,-37,-41,-13,-3,7,-24,-25,28,-9,3,5,8,-23,-8,-66,17,40,-2,-7,7,25,-17,0,35,-48,-8,-75,-1,30,4,0,-75,-8,11,-2,-12,-45,-11,20,-11,26,-82,-7,-2,1,4,5,16,-8,-4,18,27,-37,34,31,-10,22,-31,-11,-62,-104,16,23,-40,-22,22,-1,2,-28,-18,-20,-45,-35,2,19,-9,-11,-12,-26,-4,-65,9,-27,11,14,7,-60,-1,-8,-12,18,6,6,-6,-9,-40,8,20,4,7,-6,-2,-8,0,8,-14,-62,-15,0,-16,27,-4,-18,10,-9,16,-8,-7,-33,-73,8,14,-19,7,33,4,34,4,-12,-6,23,7,13,10,3,4,6,2,27,-2,0,6,30,12,-5,38,23,2,10,-50,-8,-17,-37,-80,-13,-2,-4,11,-31,15,7,19},
{34,-13,-6,-44,-16,-22,-21,-37,24,-30,-3,-96,2,6,-55,7,1,-14,-54,-5,6,2,2,17,23,5,17,0,20,-6,-2,-1,19,-22,25,44,-6,0,-35,-24,-3,-7,13,-11,-34,17,-10,-2,1,21,-17,-18,-34,42,18,8,-33,5,21,-42,22,-32,-25,7,-14,4,58,2,0,-21,-6,10,-17,0,59,-39,0,19,-10,-54,3,-7,-7,2,8,-1,-26,-12,28,40,-11,-3,2,0,0,-81,-6,-51,-83,-4,103,-8,-19,-16,2,-3,-39,-8,-36,-22,-37,2,11,-21,2,11,-24,-3,-137,6,-20,-9,11,-109,-23,-10,5,-11,23,-7,-8,-4,-10,-5,9,15,10,-11,-3,-7,-5,7,18,-20,-74,-14,40,-9,-15,-7,-57,-8,-2,25,-12,-3,-18,-67,11,3,-36,7,30,-1,37,-7,62,-7,8,6,7,24,-7,3,7,31,30,-21,6,14,28,21,4,33,15,9,8,-50,-18,-21,10,-70,1,7,-4,23,-57,-5,4,59},
{5,-10,8,-29,14,-9,-7,-30,22,-7,2,-212,-16,4,-44,0,3,-14,-7,-3,0,4,-7,19,9,-6,-22,-8,-4,7,0,-7,14,-50,11,60,0,11,-17,-14,-25,0,18,-14,-29,9,2,-10,-7,4,4,-15,2,21,-12,-6,-37,4,15,-31,15,34,4,16,-31,10,47,10,0,-3,-12,-7,-10,0,70,-29,-16,10,-14,-22,5,9,-25,43,9,0,-35,0,8,36,-19,-30,-18,-2,15,-69,-3,-63,-46,-3,104,-8,0,0,3,-7,-20,13,-37,-1,-27,-5,7,-19,-5,37,-7,34,-115,4,-12,-45,11,-88,4,-10,31,4,20,6,0,-2,-4,21,-25,24,-4,5,-4,5,2,-39,20,-12,-33,-40,34,-2,-43,1,-12,12,-1,21,1,-9,8,-60,9,9,-7,-4,26,-3,16,-2,72,-8,-67,27,21,15,-10,-6,8,10,43,4,4,6,0,11,6,12,7,-11,26,-55,-16,-13,2,-56,10,15,-2,-13,-84,4,-6,88},
{-35,-58,-8,-19,11,5,2,-15,-17,9,-7,-231,-18,-28,-27,39,4,-10,13,3,5,3,-6,7,-3,-20,-43,-6,-56,-24,-9,-22,24,-22,-14,39,2,6,-10,13,-26,0,36,-23,0,13,2,-3,-6,-20,0,26,37,-23,-26,-6,-13,3,-2,-6,-23,54,39,23,-65,6,27,18,-13,-15,-18,-9,0,-1,26,5,-15,-8,-2,-13,-5,16,-7,85,0,40,-22,-5,-18,58,-27,-81,-14,-6,19,9,-13,-47,-46,-2,33,-3,6,-20,6,-1,-8,68,-39,-12,-19,-3,-8,-2,-3,-6,23,69,23,5,2,-30,16,-48,-2,0,40,25,-26,-1,-3,-16,2,11,-45,12,-35,-5,1,5,4,-77,-5,8,7,-4,-18,3,-40,52,28,49,-7,16,6,-4,34,-23,19,-8,21,8,13,-7,-13,3,28,-3,-63,22,17,0,-12,-1,-1,-34,20,27,4,-6,12,26,3,43,11,-30,21,-35,-22,-8,-5,-52,-16,-11,-6,-61,-49,37,-4,77},
{-39,-27,3,-12,12,-5,-3,-5,-24,-35,-3,-141,-7,-39,-32,51,1,16,22,5,-2,-3,7,5,0,-11,-9,5,-50,-33,-5,-16,62,4,0,0,31,4,-10,30,5,7,29,-27,17,20,4,-2,3,-7,-14,25,46,-15,-2,-14,-2,8,18,26,3,3,35,7,-70,-7,0,17,7,-24,-22,12,-18,0,-52,9,-17,-1,14,-6,5,0,16,51,-19,54,-10,6,-15,54,1,-74,-14,-1,16,4,-14,-35,-61,-5,-51,-14,5,-7,-7,4,26,60,-28,3,-23,0,-55,-6,2,-29,9,45,115,-13,10,-9,8,-51,-13,5,37,24,1,7,-7,-37,0,12,-34,-6,-13,-1,0,4,-4,-29,-25,20,10,27,-15,-9,-10,66,21,56,-4,11,-13,0,39,-29,3,-19,-12,-8,-12,-1,-13,-7,62,1,-18,19,-4,0,-30,0,-4,-2,12,24,-1,-1,-7,52,-8,-8,8,-24,-21,-41,-10,8,3,-1,-10,-23,-1,-36,-25,4,-8,-1},
{-35,49,0,5,7,44,-2,11,-12,-46,-5,-42,-2,6,-2,25,-5,11,-32,0,6,-8,-4,-4,-5,0,18,-3,4,-21,-6,13,31,15,12,-29,17,5,13,48,9,2,-15,-25,8,-18,0,-4,-1,-14,24,-3,54,-23,8,13,17,-3,-5,25,31,-27,56,41,-13,-3,10,3,-9,1,-30,13,-16,-2,-56,-33,-16,-9,22,15,6,-1,50,14,-38,18,-26,-2,-28,3,2,-70,-16,-2,9,16,0,-29,-45,11,-81,-19,-29,-26,-1,10,7,-84,9,28,17,0,-31,-21,0,-31,-13,-81,95,-22,0,-24,10,-40,-14,1,17,17,22,7,-11,-74,3,12,0,0,17,-5,2,-9,5,-21,-48,21,-11,35,-4,8,0,-49,15,48,5,20,33,0,-13,-28,-16,10,-81,8,-25,5,27,-1,31,40,-4,23,20,-14,-12,-8,2,-19,-16,-51,6,-11,-20,46,2,-51,36,11,-11,-33,-11,20,-3,37,-6,-17,-10,28,5,-57,-9,-34},
{-16,49,-4,20,-31,20,8,-12,-4,20,1,5,0,38,16,-20,6,34,-48,-3,-6,3,3,-2,-4,-5,-16,2,41,-7,-5,-18,-4,7,24,-40,21,17,5,-6,28,-2,-74,-31,-14,-6,-12,0,-2,-2,37,-12,13,-26,12,8,24,9,-31,-1,20,-6,7,70,3,16,28,-32,-23,3,-47,17,25,-10,-25,-63,-12,4,42,43,-5,0,20,-13,-36,-7,15,-5,-19,-7,-10,-83,5,1,-1,38,-1,-23,9,26,-35,-18,-2,-105,-1,-1,6,-72,21,55,26,10,-27,-33,0,-27,-40,-132,29,16,12,-13,-6,-40,-10,-7,19,-39,-6,-5,2,-39,6,18,-1,4,22,1,-3,1,-8,-3,-23,-18,-6,-20,26,7,11,-69,-2,25,0,34,27,2,-53,0,-33,27,-15,-1,-37,8,63,-2,-66,12,25,-31,23,-3,-27,6,-4,-1,-14,-50,-3,2,-7,55,-7,-74,48,44,2,-3,-22,9,0,34,5,-30,2,66,-50,-48,4,-57},
{-11,62,5,14,-71,-11,-19,-28,0,54,-11,29,10,6,25,-69,1,34,-2,-2,5,-1,10,18,-4,-13,-5,-7,7,13,-7,-70,4,-11,34,-43,44,13,9,-44,14,3,-59,-24,2,-3,0,-9,-3,17,-20,5,-12,-8,-12,0,16,0,-7,-55,15,-31,-20,51,9,0,23,1,-10,-14,-1,32,27,0,2,-17,2,15,62,39,2,0,6,-5,-26,-30,38,6,-10,-12,-21,-30,31,5,-13,48,11,-5,15,-17,-21,-34,47,-178,-4,-3,-2,-33,27,47,32,-6,-12,-28,4,-15,-77,-80,10,28,13,1,-5,-1,-3,-3,0,-51,7,2,8,-2,-7,-28,-11,-49,17,8,4,-2,-6,23,-24,-90,12,-58,33,0,21,-15,-11,34,-9,22,-17,-2,-31,25,-89,16,49,6,-30,8,52,-5,-118,-29,36,-74,11,5,-26,5,-5,14,6,38,5,-11,-25,56,-5,-67,47,3,17,-19,-30,14,1,5,11,-29,12,51,-117,27,-3,-30},
{12,53,2,-25,-78,0,1,1,-30,50,2,29,22,-27,37,-91,-4,17,17,0,-1,-1,-4,23,-21,-22,0,-10,-6,20,-8,-85,0,-11,19,-41,35,20,50,-27,-27,1,-55,-32,25,-20,24,4,-7,13,-69,13,-2,-16,-26,-19,8,7,8,-68,0,-29,-9,37,16,1,0,66,-7,-8,0,21,19,-12,-36,-15,10,25,49,6,2,-6,35,11,-11,-25,16,-7,-20,-13,-26,39,50,5,40,36,-9,12,3,-76,-2,-39,43,-279,7,-4,5,0,28,42,28,2,5,14,-9,-26,-97,18,19,38,0,-24,1,16,-5,5,21,-38,1,3,1,27,8,-87,17,-96,8,-3,-3,-3,-8,5,-41,-49,27,-43,23,-5,32,-54,-14,15,-4,19,-49,8,-15,19,-155,-1,30,0,-7,-8,37,-7,-81,-31,31,-70,-30,-14,-20,-5,-3,-16,23,52,5,-17,-56,49,-4,-53,23,-85,-4,-24,-30,8,-17,-3,-1,4,7,8,-95,11,0,-15},
{-5,-6,8,-55,-47,12,9,3,-33,31,11,17,19,-14,29,-75,-3,0,16,3,7,-4,-2,45,-23,-30,0,0,-3,23,5,7,11,-11,10,-21,30,21,55,21,-31,0,-70,-34,43,-40,2,-3,4,14,-109,1,-9,-10,-27,-23,8,-6,-5,-54,-28,-80,-15,31,5,-20,-14,41,14,-17,-10,16,16,2,-55,-19,-55,28,5,-14,-8,-30,39,31,-5,-8,20,-1,-32,-14,-23,65,79,-2,32,4,-7,19,1,-120,5,-41,40,-335,0,-7,17,60,27,36,10,-8,7,30,6,-21,-118,143,0,28,-4,-29,-2,4,-1,-3,44,-62,4,7,-2,28,2,-97,23,-68,-3,-1,-6,-3,4,5,-55,-18,25,-43,24,3,18,-78,-33,21,-7,5,-34,2,9,30,-140,-22,3,0,-6,5,8,-6,-38,-59,24,-12,-47,-47,-12,-3,4,-20,6,10,-7,-33,-38,42,-5,-16,5,-85,-20,10,-17,19,-18,-6,-6,16,-11,-25,-47,-17,1,1},
{-38,-37,-4,-51,-6,4,-14,16,-37,13,0,16,2,-24,24,-51,-5,-6,0,-3,2,-6,2,24,-27,-52,-21,5,-11,40,-5,65,3,-6,-16,-15,14,11,34,1,-21,-6,-56,-57,35,-30,6,3,6,-8,-77,4,-25,-6,-43,-23,19,7,-35,-27,-50,-36,14,-6,4,-25,-13,5,14,-19,3,3,11,-7,-101,-5,-117,43,-23,-30,0,-27,15,33,0,4,14,-4,-13,-1,-13,61,55,0,31,-60,-13,-4,2,-114,2,-42,14,-276,-7,0,3,21,-33,-4,2,7,1,38,-2,-7,-93,116,4,12,4,-35,-18,7,-14,-7,33,-38,1,5,-1,59,-7,-101,20,-54,-5,-8,-6,6,-4,8,-61,-23,18,-4,3,-10,14,-59,-29,13,6,-9,-28,-5,31,14,-23,-28,-30,1,1,4,-4,-2,-18,-53,18,-8,-32,-60,21,0,7,-51,1,-22,-1,-24,-29,28,-1,11,-8,-107,-31,47,-20,20,-17,-10,5,29,-9,-20,-41,-41,3,5},
{-18,-10,-1,-19,-127,-1,-12,-1,-31,-9,2,14,-54,-58,5,-20,-8,-10,-10,9,-3,-9,3,0,-18,-136,-12,-6,-22,25,4,18,0,5,-7,-26,-8,-11,-15,-12,-8,-6,-30,-33,-4,7,3,-2,-3,-4,-81,-8,-169,24,-6,-6,-14,-4,-30,-51,-39,51,0,-4,6,-28,-28,-8,-3,-2,11,5,7,-7,-50,-73,-90,15,-21,16,-3,0,-6,-48,-24,1,15,3,3,-14,-8,-3,13,-11,46,-61,-12,-14,15,-111,4,-7,-12,-183,-9,1,-2,-21,-270,4,2,-3,12,18,-8,-8,-20,-10,-9,-18,-8,-31,-7,4,-13,0,3,-47,-4,1,3,-155,-3,16,10,-80,-23,-7,-5,-3,0,-34,-43,-37,-13,-45,2,1,-39,-94,-2,-13,5,-25,-42,2,12,0,-77,8,-15,8,-5,-8,-8,5,0,-20,14,0,0,-69,6,-7,5,-11,-3,-49,-10,-4,-33,28,5,-1,-69,-53,-10,45,-6,-89,-9,-1,-22,2,-6,6,-34,-47,4,4},
{-20,11,-9,-6,-3,4,-7,8,-13,-16,8,-20,-53,-6,-42,-48,-2,-25,-52,8,0,-2,-2,-7,-21,-15,-26,-3,21,44,-7,-11,-11,-18,-7,-18,-5,-62,-269,-24,-19,-9,15,-4,-21,-1,-15,4,4,-12,-1,-20,-79,8,-9,-15,1,-6,-9,-3,-53,41,-106,-20,-12,-19,26,-5,0,-19,-17,-16,-10,6,27,-8,9,0,-3,-18,-5,19,-22,-430,-88,0,11,-6,0,-14,-65,81,-47,6,0,-1,-16,7,19,9,-21,-6,-11,5,1,1,-7,-169,2,-32,12,-9,-5,-4,-4,-23,8,3,-75,-24,-33,1,-2,5,-31,-9,-22,20,-15,-3,-6,-583,-8,0,1,9,12,3,6,-4,-8,-4,3,-3,-30,-31,-6,-17,-1303,10,-29,-17,5,-68,-23,6,-9,-25,2,-8,4,-6,1,-2,-17,-6,7,-15,-44,-37,8,-32,35,0,-1,-60,-51,5,-8,3,-6,4,1,26,-39,7,15,33,4,-741,20,-17,-14,11,4,20,-13,12,-2,-26},
{-2,-19,0,1,0,0,-17,-77,13,-14,-4,32,13,-3,-83,-5,-24,-40,-68,-5,-8,7,-7,15,2,-9,-33,-5,30,58,7,-7,-10,-3,29,15,-53,-53,-45,-18,-20,-2,15,0,-1,4,5,6,4,-10,6,16,-135,24,-4,-3,-8,-7,-7,-6,-32,23,-102,-35,-37,-4,28,1,7,-22,-39,-27,-9,1,36,-9,22,-18,-6,-43,8,28,2,27,-48,8,11,-11,0,20,-36,53,-32,-2,1,8,-5,-33,0,-5,21,-16,-24,-1,-6,0,-38,-30,-5,-42,0,-11,-4,0,0,6,50,13,-38,-25,-8,-9,-10,4,-67,2,-27,11,0,3,-8,-14,5,-97,29,34,30,-7,-2,-1,-5,-5,17,-35,-56,-25,-9,-14,65,14,-38,-48,6,0,-26,-13,-9,-60,11,-16,-17,1,27,4,15,-1,-35,-4,29,-50,19,15,56,6,-9,19,-10,2,-3,9,6,-2,0,49,13,10,25,-21,-6,6,-31,-52,-10,3,-3,3,-3,1,5,25},
{1,-16,8,-9,-36,-6,-26,-56,30,-12,0,87,0,7,-84,-7,-11,-15,-67,-7,-1,-8,-9,27,16,-11,-18,-5,34,-13,2,-8,15,-5,46,33,-31,-26,-51,-5,-3,2,3,-5,-23,19,0,-3,0,26,-6,-12,-91,37,8,-2,-12,4,7,-15,-9,-63,-79,-29,-25,4,42,-1,-20,-16,-15,10,-19,0,13,-9,15,-4,-6,-34,-3,13,0,25,3,1,10,-3,4,5,-31,-2,-22,-6,13,-15,6,-31,-110,13,69,-8,-19,2,-6,-3,-44,-20,-15,-39,-1,6,9,3,-2,10,27,11,-21,13,-10,4,-5,-35,-33,4,4,-1,6,6,6,-7,-10,-53,33,23,22,-2,3,-7,-2,7,21,-14,-135,-5,17,-10,49,6,-55,-46,0,14,-33,-5,-26,-40,14,5,-35,-8,43,-7,20,6,36,-9,40,-37,-3,33,8,3,8,56,-4,-15,-9,14,3,7,0,84,19,23,17,-7,-18,-22,25,-67,-6,19,3,2,-10,-1,-10,44},
{5,0,-4,-25,1,-11,-33,-56,22,0,8,-24,4,11,-76,-18,-7,-5,-54,-5,-4,-11,-2,45,30,-14,3,2,29,-53,7,0,-13,-51,49,67,-39,-18,-49,-6,-16,3,0,-9,-30,17,-7,-8,5,24,-2,-17,-55,25,1,-2,-22,-3,15,-31,9,-78,-63,-23,-5,5,57,0,-22,-7,2,21,-19,-8,55,-27,5,14,-23,-5,-8,18,-4,30,4,-3,-16,-12,7,10,-15,-46,-15,-11,17,-35,5,-21,-72,11,120,-7,-6,-5,7,0,-40,-7,-32,-16,-8,1,13,-8,-6,9,21,19,-35,6,-9,-9,13,-104,-8,-10,11,-2,15,-2,2,-8,6,6,31,5,35,3,-7,0,3,-2,33,-20,-131,-11,20,-8,11,-9,-57,-37,-5,33,-34,-9,-21,-17,9,5,-41,-4,32,0,16,-2,58,1,-28,6,5,27,-46,4,-1,77,-9,-8,0,22,-2,9,-1,107,23,4,0,-35,1,-27,56,-51,-2,26,-11,7,-22,-2,-9,74},
{-9,-19,0,-1,27,18,-20,-34,13,4,-2,-191,-1,-21,-36,3,-1,0,-5,0,-8,-13,-3,19,-1,-19,-13,2,3,-114,4,-11,5,-77,9,41,-49,-20,-21,20,-29,-9,33,2,-32,25,12,-9,-7,13,14,2,-13,2,-10,-3,-4,-3,6,-19,11,-46,-39,-1,-22,19,48,31,-25,5,-3,3,15,8,31,6,-15,9,-15,-11,-8,16,-7,99,8,20,-33,-4,-19,17,-14,-70,-10,-4,49,-10,-11,1,-44,0,72,-12,9,-11,-1,3,-27,30,-26,-11,4,-15,9,12,0,-5,70,61,-21,23,0,-13,19,-33,4,4,10,19,2,-7,4,-6,3,35,8,-1,9,8,8,0,-4,-50,16,-10,-71,-21,11,-1,-8,27,8,-19,-10,21,1,2,-2,3,21,8,-11,-1,28,7,-11,8,29,-8,-124,33,43,15,-35,7,4,4,-6,28,9,14,-3,-16,7,73,13,-20,10,-53,0,-9,40,-54,6,12,2,-32,-28,25,3,73},
{-35,-37,-7,18,-4,28,-6,-12,-7,5,0,-164,-8,-21,-2,8,-2,16,18,-8,3,-5,6,2,-31,-4,-10,-4,-16,-98,-5,-7,34,-29,-5,-21,-25,1,-21,28,0,-9,40,3,-8,14,11,-1,1,7,23,34,0,5,-14,1,39,4,-10,8,-22,-22,-10,-27,-12,24,9,18,-2,10,-8,29,9,-4,5,28,-27,2,4,-4,8,5,-11,65,-16,-1,-16,-11,-20,20,7,-52,-4,13,9,0,-1,13,-44,19,0,-30,18,-10,4,2,26,48,-17,-21,4,-5,-4,15,6,-34,37,61,-5,10,26,15,0,-1,-17,-3,-6,37,0,3,-6,14,4,33,28,3,0,-12,-3,0,3,-41,-17,6,6,0,3,8,12,57,36,-12,-4,15,-2,-2,-33,19,6,0,21,-3,5,-6,-13,7,65,-9,-86,22,12,-14,-72,8,6,-46,-28,34,-1,26,-13,-46,11,56,24,-16,-19,-50,15,20,15,-24,-8,8,-2,-21,-1,26,-9,24},
{-4,-14,-9,2,5,47,-3,-10,-8,-7,-6,-39,26,4,8,16,7,17,-13,-1,-5,-9,3,-9,-20,11,7,0,13,-51,-5,0,46,-4,15,-43,-20,14,-18,18,44,-6,46,-6,20,-3,10,-4,8,9,9,7,-5,0,-5,8,40,4,0,-4,-19,-30,29,-36,-8,15,-2,11,0,5,2,19,-14,-4,-36,-10,-12,16,0,-2,-5,-2,41,9,-29,-25,-33,-9,-8,12,10,-34,-4,0,-1,15,17,26,-24,32,-85,-41,-2,-6,-3,-9,31,-68,-9,-33,3,1,-14,22,5,-36,-2,-24,19,7,11,2,-16,19,-16,0,-19,55,25,-5,-6,-3,-3,18,33,8,16,-11,2,8,4,0,-19,35,5,-11,11,-5,28,19,31,-14,7,36,21,-3,-68,16,13,-5,0,0,-16,-6,3,-8,40,16,-47,17,0,-19,-25,-1,5,-46,-42,17,5,38,-12,-62,-3,41,11,1,-28,-51,15,48,-9,22,0,-21,-12,47,29,-33,-6,-29},
{-1,33,-3,7,10,33,-1,-18,21,-4,-1,85,51,28,7,9,11,14,-40,-2,-1,-8,-7,-32,-4,6,23,2,64,-38,5,-10,3,31,51,-41,-29,35,14,19,43,-5,-48,3,17,-17,-19,10,0,12,42,-34,9,-13,10,31,18,1,21,-35,0,-55,28,18,1,3,-4,12,7,0,4,6,-11,-5,-44,-21,-2,8,-3,7,-4,3,34,-51,-42,-29,-41,-2,0,15,28,-6,-2,-10,10,18,10,48,-51,24,-58,-30,-18,-17,0,6,5,-104,-1,-9,-14,3,-5,-9,10,-39,-16,-75,-13,7,11,0,17,12,11,2,-15,-21,23,0,-2,-13,-1,23,23,13,21,-7,-6,4,-4,6,9,-1,-29,-15,1,0,2,-48,40,-14,6,39,47,8,-71,10,13,32,-32,-8,-12,4,42,-8,-14,33,-27,-20,9,3,10,-5,-8,-19,-37,-56,-4,11,10,-24,-5,2,9,42,12,-12,5,68,4,32,-9,-40,-1,70,15,-8,8,-71},
{-31,16,0,21,-18,-28,-6,-45,64,31,1,25,26,22,35,-30,7,44,-3,-3,0,-8,0,-13,28,-13,25,0,42,-14,1,-51,-25,49,54,-63,0,43,-4,13,47,2,-51,8,12,-15,-40,6,7,17,3,-42,21,-16,-6,51,31,4,-37,-58,-19,22,-5,56,12,0,1,-47,-1,7,-6,23,-2,0,-30,-6,10,-16,-1,32,-5,0,-32,-48,-29,-31,2,6,19,23,11,18,-7,0,0,10,2,12,-8,16,52,3,12,-29,-1,3,1,1,2,69,-7,-9,-5,-67,1,-38,-20,-17,-32,10,20,-5,9,-34,13,6,5,-65,13,-5,6,-11,7,37,-5,-36,17,-1,-4,6,-4,-10,5,-53,-27,0,8,7,-29,15,29,0,0,16,-26,-2,-47,35,-7,20,12,4,-20,-8,80,3,-43,34,21,0,28,28,-4,7,-7,45,-40,-54,-1,-18,15,54,1,12,10,2,2,4,-3,87,17,-6,-2,-28,0,38,-52,10,1,-25},
{1,39,-8,12,-24,-41,-8,-48,45,42,3,-4,8,0,32,-72,4,32,-19,-4,8,-9,0,25,3,-40,14,-7,22,-19,9,-94,-27,-2,38,-53,44,16,-16,-11,14,0,-7,18,-12,-13,-2,0,0,25,-34,-3,-3,-19,-3,19,63,-6,-29,-38,-35,-7,-2,66,29,12,13,-3,-6,0,0,24,10,-10,4,6,51,8,14,30,-2,-19,-42,-41,-20,-52,55,3,-6,0,6,29,-12,-2,24,50,-6,5,13,4,27,3,39,-73,2,1,-11,-55,3,68,3,9,4,-33,-2,-36,-20,-7,29,26,10,9,-9,29,-15,7,-11,-10,11,3,-1,15,10,-12,-2,-73,42,-8,-5,-5,-4,45,-6,-31,-34,-5,15,8,37,22,17,-8,0,-13,-61,-1,13,43,-61,0,0,2,-41,-3,64,1,-76,-4,35,-37,16,2,-29,1,7,47,-38,14,7,-33,-6,88,2,20,3,-60,-3,-51,6,32,3,-36,-2,45,-10,29,-55,30,0,32},
{16,49,5,-3,-52,1,14,-10,16,66,-2,15,34,-14,40,-92,1,0,-18,8,9,-11,11,57,-8,-47,20,0,33,-49,-8,-68,-27,-26,26,-32,33,-1,22,-33,-53,7,-18,18,-8,-47,27,-2,-7,11,-61,10,3,-30,-8,0,31,3,8,-16,-47,-54,-52,34,12,1,13,49,-26,1,3,4,5,-12,44,22,50,43,-7,-4,4,-18,-4,9,-26,-80,44,-10,-44,-13,-18,22,7,-3,44,35,-10,6,4,-27,19,-7,37,-71,7,-3,-9,-55,3,17,11,-2,17,56,5,-28,-24,27,73,31,13,1,11,63,-19,0,42,-31,21,4,-5,43,8,-76,27,-41,28,10,0,4,6,12,-23,-55,-10,-46,19,-2,33,-9,6,-14,0,-36,-65,14,23,45,-82,-15,28,3,-14,3,22,-4,-60,-24,19,-62,-39,-23,5,-6,7,-33,-9,35,3,-25,-14,84,2,44,-33,-108,5,-18,15,12,-9,-14,-1,62,2,0,-9,32,-3,0},
{37,-4,-8,-24,-68,19,6,9,37,81,-4,15,24,-9,46,-80,-8,-13,4,-6,0,1,-8,57,-23,-31,20,3,21,-38,0,46,-9,-18,2,-26,10,12,36,-5,-67,6,-20,7,19,-75,-18,2,-4,7,-91,-28,7,-13,-25,0,-3,-6,-3,-29,-104,-111,-44,16,14,-28,-9,50,-6,-12,-11,11,-6,4,2,6,-35,49,-61,-15,7,-34,21,18,-12,-57,31,-4,-55,-6,-27,11,60,-7,32,7,6,-7,4,-43,18,-31,12,-30,3,-7,-5,20,6,22,12,0,-6,57,-2,-26,-33,121,34,22,7,-31,21,35,-15,2,64,-55,41,1,0,23,-2,-47,36,12,12,7,-5,1,-8,-5,-31,-54,21,-50,14,4,12,-24,-28,-14,2,-56,-33,15,38,52,-77,-17,12,-3,-5,-5,8,-7,-42,-59,6,-16,-60,-48,17,3,8,-37,-4,5,6,-64,2,64,3,52,-25,-118,-12,23,-8,21,2,-5,-5,52,-1,-31,17,-3,-2,10},
{0,-36,0,-45,-43,4,4,12,-36,40,1,-1,24,-19,32,-27,4,-11,-7,1,3,3,-6,38,-25,-22,-3,-8,-9,-1,0,84,8,-17,-8,-37,-6,20,28,10,-40,4,-24,-18,18,-30,-11,-3,-6,-9,-68,-24,3,-2,-18,-19,6,4,-27,-26,-33,-64,9,-6,4,-37,-30,9,24,-12,7,5,18,-7,-106,-14,-138,52,-64,-14,-5,-44,2,14,4,-3,13,-1,-10,10,-23,19,38,4,32,-19,-5,-1,0,-74,15,-40,3,-242,1,-9,-3,37,-38,11,-4,8,-16,34,-5,-15,-41,192,14,11,4,-13,-7,19,-3,-7,41,-40,7,-1,-8,41,-6,-73,24,50,3,-1,-3,0,5,9,-46,-13,-2,-4,1,0,7,-66,-34,-22,-7,-65,-3,8,22,27,23,-42,-12,-4,8,4,-3,-8,-40,-32,6,-7,-34,-75,53,2,4,-36,-6,-34,-7,-36,-19,23,0,23,-39,-46,-32,42,-6,37,0,-5,-1,39,4,-11,-13,-41,0,15},
{-16,-22,-2,-44,-13,-1,-8,2,-48,-26,9,-11,-4,-32,29,2,5,-4,6,0,0,-5,-8,-5,-18,-49,-18,-6,-18,-6,-2,28,-9,-9,-18,-2,-19,0,-22,-18,-13,-6,-6,0,-3,7,-44,3,0,2,-65,-23,38,10,-19,-29,-38,4,-14,0,-70,23,10,-18,9,-17,-54,-15,-9,2,10,2,15,-5,-70,-24,-297,-27,-21,7,-2,-32,-12,43,8,0,4,3,-9,-6,1,12,8,8,32,-75,-14,-24,5,-93,11,-18,1,-24,0,-5,-16,10,-153,17,8,6,-6,32,-10,-16,10,52,-9,-12,3,-26,-26,13,-10,-5,15,-21,14,0,-4,63,-9,-60,6,-32,-45,-7,-6,-5,-4,-9,-21,-21,-16,-29,15,-13,3,-18,3,-54,-10,-40,-46,-17,18,26,42,-11,-18,-6,-2,7,0,-5,-61,-9,-14,-1,-10,-12,33,-6,-5,-35,16,-31,2,-15,-14,-10,-3,15,-82,-73,-22,59,2,-9,5,-14,-14,7,-7,0,-13,-21,0,-2},
{-14,19,-7,-4,-49,-3,-11,-4,-8,2,-3,-4,6,-28,-70,-7,-16,-11,-70,-4,-6,6,6,-6,-40,-7,0,-2,18,26,-7,9,-28,0,4,-47,4,-102,-255,-5,-53,8,31,5,-8,3,1,2,1,12,-10,-21,-114,0,-7,-33,-2,2,-9,-3,10,46,-110,3,-10,-3,41,1,3,-19,-10,-10,-21,-4,53,-42,4,-24,3,-14,1,20,1,-18,-688,-24,12,-2,5,-35,-96,59,-40,-10,1,1,-6,11,30,0,16,0,-2,-5,-5,-4,-10,-121,25,-20,-12,-4,-9,-2,3,-4,-35,1,-47,-17,-11,4,-2,6,-27,-8,-34,17,-1,5,6,-461,-8,-55,30,-4,30,3,6,-4,6,-1,2,-2,-25,-46,0,-14,1,-3,-4,-29,4,-41,-114,-10,31,-38,-1,0,8,-3,-27,8,0,-4,-27,-26,-7,-49,-8,-7,24,5,1,-5,-31,1,-6,3,-9,-49,7,-11,-37,-12,4,58,3,35,1,-12,-19,32,-7,22,-5,0,-9,14},
{0,-18,1,0,-26,9,-10,-101,-2,-3,8,81,0,4,-96,-18,-5,-22,-66,2,1,-7,0,21,-8,-9,-17,4,40,63,-9,-20,44,1,66,41,-88,-64,-47,-12,-33,0,12,6,-4,6,8,-7,-6,0,0,9,-131,25,5,-16,-14,-4,-15,-8,-2,2,-72,-93,-17,9,33,5,-8,-13,-12,-11,-3,1,43,-10,9,-38,-28,-26,4,19,0,46,-38,5,10,-9,-7,-18,-55,-1,-31,-10,1,6,1,-70,28,5,29,-7,-4,13,0,0,-41,-21,-2,-16,11,2,-3,24,-3,5,36,13,-21,1,-7,4,2,23,-34,5,-43,4,9,6,-4,-8,-1,-77,45,18,34,-5,-7,5,6,7,15,-39,-123,-16,-4,-8,56,0,-43,-69,3,-19,-34,-17,13,-36,3,-3,-23,-8,22,0,-8,0,32,-21,42,-8,25,12,41,-5,-5,15,-20,-13,0,7,2,-2,3,60,-6,12,37,24,7,-19,43,-42,-12,12,-7,5,-3,-2,-4,26},
{6,17,8,-6,-29,-6,-34,-64,21,0,-8,160,0,11,-84,-16,-7,-1,-79,8,-1,-11,-3,24,17,-15,-15,7,32,-7,-4,-8,39,-4,52,20,-34,-21,-74,4,-15,6,7,-3,-2,16,0,-1,-10,26,-3,-37,-73,18,-11,-4,-7,0,-7,-19,9,-119,-69,-57,-16,5,35,24,-32,-4,-1,16,-8,-4,59,-8,24,-7,-38,-17,6,24,8,25,-3,-17,13,0,5,-30,-28,-30,-43,-10,11,-21,-2,-51,-109,3,85,3,-18,-5,3,4,-46,-17,-14,-18,22,-3,9,13,3,3,39,11,-17,13,-4,-7,12,-47,-17,0,-4,-3,13,0,5,20,-6,-49,36,12,45,-5,-2,-4,-4,41,18,-23,-175,1,13,-11,47,-2,-56,-120,1,-1,-55,-13,-2,-23,9,7,-48,6,29,4,14,-8,74,-19,20,-33,8,23,-6,7,-2,57,-12,-10,-3,17,3,-10,2,81,2,10,7,11,3,-24,62,-29,-2,21,4,17,-9,-6,2,55},
{5,11,8,-2,-4,0,-5,-55,28,-8,-7,109,3,-3,-43,-32,-14,7,-44,0,4,-6,5,20,27,-26,-14,11,20,-61,6,-3,40,-52,34,30,-37,-19,-43,9,-40,0,21,2,-17,10,-2,-7,-4,23,2,-24,-22,-15,0,0,-6,4,-25,-20,43,-114,-61,-27,-7,13,59,18,-27,4,11,7,-6,5,53,-15,6,9,-33,2,0,15,-1,41,-2,-9,-6,-12,0,-18,-15,-99,-45,-4,59,-39,13,-36,-62,11,56,13,1,-10,5,1,-36,17,-16,-21,19,-8,14,0,0,-3,83,54,-4,24,-1,-10,25,-22,7,-6,-6,4,16,1,-8,23,0,15,31,-9,57,-8,-4,2,1,-1,26,-26,-169,-34,30,-5,24,20,-14,-85,-8,16,-41,-3,-8,10,9,26,-54,5,26,-8,-4,8,62,-12,-51,-32,25,17,-32,-8,1,42,-27,0,-9,5,0,-19,2,94,2,-17,-23,16,2,-19,70,-32,3,28,13,12,-33,6,2,37},
{-19,-31,-1,29,9,39,7,-13,3,-13,-3,-85,-8,-34,8,-13,-15,20,0,2,0,3,5,4,-31,-12,-28,2,-9,-101,-5,-16,20,-62,-17,-28,-24,-4,0,35,-38,6,32,10,-19,7,3,-9,1,8,27,-1,31,10,0,18,13,0,-10,1,19,-62,-27,-15,-9,21,30,11,-14,20,19,16,23,3,26,24,-21,19,-8,17,-4,2,-20,91,0,-1,-29,-10,-7,-11,-25,-117,-37,0,8,-20,-3,-5,-34,13,14,-15,11,-6,6,-1,15,55,-8,-17,40,2,0,2,-6,-28,86,104,3,17,16,5,29,11,4,0,-29,18,10,1,-6,27,3,30,42,-21,28,-7,4,-5,8,-64,7,-24,-67,-28,-1,6,-10,28,30,-65,5,-5,-10,-2,-14,28,5,22,-11,6,25,0,-47,-7,17,-9,-109,-24,45,-11,-47,-9,-7,-64,-24,38,0,13,0,-15,4,66,2,-22,-19,18,11,5,52,-18,0,43,-7,0,-13,13,6,33},
{-20,-72,8,41,-9,40,-3,24,-18,13,0,-112,-3,-64,32,1,0,37,32,-6,3,-2,6,-16,-45,-6,0,9,-20,-22,5,-7,31,-9,-32,-54,1,-5,5,34,7,6,20,1,-11,19,-3,-6,-2,13,1,-8,32,31,4,2,38,0,-22,20,-37,-6,-27,-18,-46,16,-17,-12,8,4,19,1,7,2,-20,43,-16,9,-21,8,3,-14,5,50,-24,2,0,-11,4,-3,-11,-73,-28,-7,-30,21,11,-28,8,-2,-75,-12,22,20,8,0,59,31,4,-31,33,0,-9,24,-1,-12,60,38,36,21,16,21,0,21,1,0,-40,29,3,-1,-10,24,-3,27,21,-18,-4,-10,-6,-5,-1,-55,-16,16,-22,-13,-2,8,17,21,13,-34,1,-29,5,-10,-23,18,1,0,17,-8,-2,-2,-18,0,49,0,-5,-10,6,-28,-33,3,-6,-50,-13,35,0,33,-13,-33,3,75,-5,0,-45,3,37,33,-15,25,-11,34,0,19,11,-6,-6,-4},
{26,10,-6,30,22,48,0,24,12,-16,3,38,34,11,5,14,8,31,-24,6,1,-3,9,-23,-10,10,-14,7,4,26,-2,20,50,9,3,-32,-7,-10,-9,6,19,-4,-28,14,5,-15,10,-1,0,22,24,-32,-6,32,10,3,30,-4,-42,9,-30,-80,-19,-21,-20,-20,-38,5,4,-10,22,-12,10,-1,-67,20,-8,23,-30,4,-6,-5,30,-55,-12,-6,35,2,19,-9,-1,5,-7,-12,-21,28,17,27,25,16,-85,0,-6,17,2,5,12,-44,-4,-61,6,8,-3,42,-2,-15,43,-106,83,-1,-4,17,14,53,-12,2,-50,13,19,8,5,-12,-5,-4,10,0,-1,-1,5,-3,8,2,-23,19,-14,29,24,-2,44,-18,-13,-29,0,-30,0,8,-21,-9,24,-20,-34,0,0,4,5,-4,18,-12,19,-8,-26,-30,-3,0,7,-1,-5,8,-3,23,-12,-41,-7,18,-10,32,-41,24,17,36,-16,19,2,13,-9,66,45,-24,8,-122},
{12,26,-6,31,17,23,-3,-9,17,-18,-3,71,54,45,-19,-5,-1,0,-49,-4,-7,-1,-8,-26,6,12,1,-10,37,43,8,0,-4,11,27,10,-41,-12,0,22,35,9,-5,2,-21,-28,6,3,-4,44,33,-50,-19,38,0,35,25,-3,-45,-46,-16,-27,-34,-28,2,-58,-35,-46,-1,17,25,-7,13,7,17,26,12,-5,-39,11,0,-6,-16,-68,-13,-29,5,0,47,28,14,0,10,-15,-11,15,0,44,5,8,34,7,-63,18,-1,1,-45,25,-5,-23,-1,2,-22,16,6,-10,67,-47,25,-30,-20,24,50,25,14,-7,-61,-53,22,3,4,-17,4,-12,21,19,5,-12,1,0,-4,-2,14,-16,-8,12,18,2,10,-12,9,-16,10,-27,-5,9,-18,9,34,2,-37,8,16,5,-4,-3,-15,14,17,-17,-2,12,17,6,0,27,9,-63,-5,6,-40,-15,-4,-1,0,22,27,83,-2,45,33,29,-11,-12,-11,50,-15,19,-1,-83},
{-44,11,4,45,-25,-50,1,-32,26,12,4,0,22,14,9,-6,3,13,14,3,0,2,-2,-12,42,-5,2,0,20,-2,4,-43,-39,14,24,-19,-12,-6,-31,-24,31,-5,21,9,-20,-9,-8,5,-7,9,-11,-61,23,2,20,63,16,2,-35,-53,31,53,-26,3,15,-17,-23,-65,8,32,33,-16,-1,5,10,23,18,6,-27,20,6,-12,-49,-41,-6,0,-24,-4,35,8,20,-4,-20,3,0,-30,-1,19,7,13,96,46,-24,-7,-4,4,-50,51,-6,38,-11,-13,3,-58,4,-32,52,42,47,-7,-11,27,33,-18,1,5,-51,-14,30,-8,0,-9,0,1,3,-7,46,2,-6,-2,-2,-26,4,-25,-45,31,38,0,-24,51,-26,-43,5,-28,-21,8,-20,17,17,-3,7,3,18,-6,22,0,-11,55,13,20,22,2,6,1,0,34,-13,-15,1,-13,-3,29,4,41,9,11,-10,31,-31,64,42,24,-4,-28,-4,16,-43,18,0,36},
{-5,25,0,5,32,-49,-8,-1,29,4,5,-25,-3,14,44,-41,-3,30,3,-1,6,0,-3,31,23,-35,6,0,41,-31,7,-118,-42,-14,-12,-22,41,0,-83,-26,-13,1,64,9,-6,-3,-1,1,0,8,-3,19,38,-2,18,41,38,2,-46,-15,83,35,9,18,16,43,-14,-35,1,11,0,-13,-4,2,31,-17,42,36,-28,32,-2,-55,-59,-25,-10,-47,39,1,-24,-13,30,-1,-42,2,34,-4,11,-1,11,24,49,35,21,-57,2,0,-26,-67,5,20,-23,-7,9,-35,2,-25,37,6,89,-2,-10,11,-26,0,-25,-6,-2,50,36,0,0,4,6,-56,5,-85,56,7,6,8,-6,44,-8,35,-65,23,2,7,13,23,-36,-37,0,-56,-30,11,13,42,1,-2,-4,-7,-17,0,28,2,-17,16,-3,-21,20,-15,-17,-1,8,5,-33,-16,9,-18,1,56,9,50,-16,1,-26,-18,-9,34,-1,-3,9,72,-13,-6,-18,-15,9,74},
{24,6,8,-6,-14,-31,-1,23,12,24,8,0,36,9,41,-50,10,8,-40,0,10,4,-4,55,-28,-25,3,0,93,-99,3,-25,-50,-30,-6,-8,27,6,-52,-54,-8,-7,37,1,-18,-47,-10,5,8,-9,-21,-12,37,4,8,-11,13,3,0,-9,-14,-83,-3,12,-4,26,-2,-7,-17,4,-21,-14,-16,-1,54,-12,10,50,-38,-6,1,-26,-40,27,-24,-83,27,-9,-65,-15,-5,-26,-9,4,18,-9,7,-31,33,17,8,4,13,-23,5,0,-12,-48,24,-26,-7,0,-2,45,0,7,38,-6,90,5,0,-5,8,49,-46,-3,27,35,20,7,-9,25,-6,-74,24,-33,28,-4,-6,7,8,45,-13,-16,-28,-27,-17,12,29,23,-34,-32,-3,-67,-76,11,67,41,-32,-13,30,-2,-16,-6,-1,8,-27,-5,-19,-62,-38,-34,-7,5,-4,-33,-1,27,1,-28,-9,58,-5,66,-30,-49,2,-11,18,2,0,-2,1,67,0,-27,22,6,-1,37},
{31,-17,-4,-14,-39,14,-10,14,37,18,11,21,18,3,21,-49,-10,-12,-14,1,-2,-1,2,58,-35,2,4,4,57,-77,-5,51,-28,-31,-6,-21,-4,13,-33,-23,-49,0,36,10,-15,-48,-25,-4,9,-12,-45,-76,24,-6,-19,-16,-22,-9,-23,-41,-79,-132,-25,-13,-15,-8,1,24,-11,-4,-29,-13,-12,11,5,-15,-76,31,-78,-11,-3,-26,7,22,-17,-86,12,-12,-44,0,-27,-49,38,0,-24,20,5,-25,34,-3,23,-18,0,16,4,-2,-12,41,3,-8,17,3,-32,45,2,15,52,33,55,-9,-9,-26,21,51,-12,6,53,-12,-1,-2,2,10,4,-30,11,47,0,8,5,0,4,16,-1,-71,-10,-42,-11,7,23,-13,-42,-45,-4,-48,-56,2,66,36,-20,-8,9,6,-9,0,-7,1,-40,-38,-20,-11,-37,-33,25,-7,8,-36,15,34,-8,-46,4,43,-5,63,-33,-55,11,43,11,4,37,15,1,32,-1,-54,40,-3,5,15},
{14,-44,-6,0,-48,10,-9,1,-1,33,3,5,23,-38,32,0,3,-9,-5,-4,4,-8,10,21,-24,1,24,1,17,-42,-3,67,-5,-10,-35,-29,-24,16,12,3,-32,2,10,7,-25,-17,-45,-7,3,5,-45,-82,12,-3,-17,-19,-14,0,-22,-19,-8,-91,-2,-2,-1,-34,-28,0,15,-4,-6,-7,-1,-9,-66,26,-214,4,-68,-16,-3,-28,0,11,13,-64,-1,0,-4,-2,-17,-39,10,-4,-4,-2,1,-11,11,-39,24,-44,0,116,3,5,-10,58,-23,-10,8,-6,-30,24,0,27,41,128,21,-23,-23,-9,-6,18,14,6,7,-41,-2,0,-5,19,-7,-42,15,148,4,4,3,0,7,-13,-10,-21,-17,-34,-1,-4,10,-47,-18,-61,-5,-52,-10,-5,16,33,28,-22,-22,-6,3,8,-5,1,-54,-39,3,18,-20,-50,56,-2,6,1,0,-18,7,-23,-8,-17,-8,38,-65,0,0,54,5,19,22,2,1,16,-5,-15,9,3,-2,8},
{1,-40,8,-40,22,-18,-2,6,-55,-29,8,-3,-34,-54,16,14,-11,-7,-15,-3,-1,-3,-6,0,-38,-12,6,-8,-11,-16,2,53,-10,-16,-27,-1,-9,6,-16,-24,-27,0,-10,-1,-11,-6,-10,-1,-3,-17,-24,-37,60,5,-13,-41,-32,-9,-10,-2,-11,36,23,-6,1,-23,-80,-24,-5,1,13,15,18,7,-80,-25,-308,-36,-17,11,0,-37,-14,52,-36,-25,8,-5,-22,-1,-11,-22,-3,-4,3,-340,-18,-2,1,-59,15,-26,14,71,0,4,-16,5,-119,33,12,-6,3,17,-7,-4,43,76,22,-17,8,-21,-35,13,0,-1,0,-13,17,3,-5,33,3,-9,5,20,-38,0,-4,0,6,-23,18,-16,-31,-24,24,-14,6,-9,13,-55,-7,-56,-25,-8,14,14,67,-13,-20,1,-14,-7,-11,-5,-42,-17,-19,10,0,-25,31,1,5,21,12,-31,4,-9,7,-92,-7,19,-106,-36,-26,52,-3,-38,4,-19,-19,6,5,4,-5,-13,0,6},
{-8,21,-7,-22,-48,-8,-7,-13,-22,-8,-8,14,-35,-36,-60,0,-12,-19,-51,0,5,3,-4,-11,-11,-9,-2,-3,0,6,5,-13,-26,6,2,-79,13,-104,-159,-2,-64,3,23,1,3,25,-1,2,2,15,-12,-7,-1166,0,-12,-31,-2,-8,-27,-3,4,-16,-211,-6,7,0,19,-8,5,-20,-6,6,-28,6,30,-41,11,-43,2,-9,0,24,10,-48,-360,16,0,-6,5,-36,-82,26,-30,0,-8,3,-9,0,31,-7,16,2,-11,2,-1,4,-11,-69,28,-13,-16,-1,3,-18,-11,-7,-36,-2,-70,-10,-16,-17,-1,0,-24,-3,-51,7,-1,6,-9,-291,2,-37,23,-7,30,-6,-5,2,-4,-10,-6,1,-22,-57,-1,-18,-52,-6,-18,-27,-6,-66,-157,-8,44,-32,0,-12,10,1,7,-8,3,0,-48,-28,-22,-31,2,-6,13,1,3,-225,-26,-21,2,0,3,-259,0,0,-47,-2,24,26,4,-429,-7,-18,1,39,-11,11,-14,-8,-6,5},
{-4,-19,2,-13,-30,-1,-20,-87,-4,5,3,91,-3,7,-65,-26,2,-16,-71,4,4,-8,-12,31,0,-7,-8,2,25,33,2,-25,46,16,81,-11,-49,-59,-43,-15,-31,1,10,7,1,4,-5,6,6,19,-3,-17,-78,28,-7,-19,5,-4,4,-6,-10,-57,-54,-76,-11,0,0,0,-25,-19,-5,1,-2,2,3,-13,11,-34,-15,-25,-1,-1,0,42,-58,-10,31,-12,-10,-26,-39,-6,-16,-12,12,3,3,-68,31,0,38,-9,-19,12,3,-3,-32,-25,11,-8,21,-11,-1,21,-9,7,25,10,-9,4,0,-2,0,-3,-37,6,-38,-1,2,0,-7,14,-5,-65,39,7,26,-7,5,-8,8,17,8,-19,-108,-4,7,4,42,-8,-24,-130,-9,-40,-54,-2,30,-21,9,0,-27,1,19,-8,6,7,19,-33,36,-21,39,5,12,0,0,39,-16,-14,-9,1,6,-17,4,39,-27,2,16,40,5,-10,52,-36,-3,28,-7,-10,-5,1,5,35},
{15,13,-3,-2,-6,-17,-22,-72,27,5,-1,185,0,22,-54,-38,-8,0,-66,-5,1,-2,-4,28,27,-13,-4,9,35,-37,6,2,81,-39,42,-18,-45,-33,-64,10,-34,-8,4,1,-20,20,-17,-2,0,24,-8,-65,-38,11,0,-2,-20,3,-10,-1,24,-126,-60,-66,-23,14,-5,5,-37,-4,-2,25,-13,-1,-9,-18,6,14,-27,1,-7,-6,1,20,-3,-24,-1,-7,4,-35,-19,-75,-38,-2,19,-21,-5,-109,-68,14,54,-5,-7,6,6,1,-30,5,-2,0,37,-5,7,29,-11,0,51,19,-4,13,4,0,25,-15,-19,-3,0,-1,6,-1,8,22,2,-15,43,-9,45,3,-8,-4,6,28,13,-13,-140,-17,11,-3,35,8,-45,-140,-5,-16,-63,-7,29,19,9,8,-53,-3,23,0,3,2,47,-19,13,1,-9,16,-26,-4,3,80,-8,-17,1,-1,4,4,-3,70,-6,-10,-18,50,-1,-13,68,17,-1,13,9,-17,-5,-3,-10,23},
{20,0,-5,-1,11,15,-12,-32,5,2,2,109,11,13,-22,-26,-9,14,-28,-4,-6,-4,11,25,6,-12,-14,1,-16,-106,-4,-8,69,-69,14,-18,-44,-27,-36,24,-32,-5,37,2,-37,3,-13,-3,-2,-7,-1,-70,7,-39,18,8,-10,6,-9,0,28,-91,-40,-60,8,26,-9,19,-17,2,19,23,4,0,-22,-1,-16,25,-19,0,0,-23,-3,66,0,51,-21,-9,-5,-8,-22,-144,-39,-8,29,-30,-8,-50,-46,22,25,-11,15,-9,7,9,-11,37,11,14,42,8,11,21,-7,-5,99,52,15,15,9,8,42,29,-17,-1,0,20,5,0,-10,17,5,10,38,-3,50,-10,7,-8,3,-9,-2,-10,-124,-29,10,-4,20,21,-13,-97,0,-3,-50,0,24,49,8,20,-41,3,8,-4,-32,-4,-21,-22,-62,39,12,3,-14,-9,0,15,-6,8,9,1,4,-7,0,87,-22,-26,-27,66,-3,-13,39,-24,-1,1,0,-35,-19,25,4,0},
{9,-81,2,17,23,43,0,-9,7,15,3,-50,-22,-43,17,-1,10,31,35,0,5,10,4,-5,-60,-15,27,-4,-30,-83,3,-18,25,-34,-23,-46,0,-4,41,15,-22,0,-5,7,-47,37,-29,-6,1,-14,7,-49,52,0,19,2,-7,-7,21,10,1,32,-2,-33,-21,24,-40,10,22,2,27,-4,0,5,-84,34,-29,9,-6,7,-6,-36,-31,106,8,51,-48,-6,10,28,-29,-114,-26,-3,-41,10,6,-27,-26,4,-42,-20,25,10,4,12,36,65,17,10,33,-4,8,14,-1,6,75,39,29,4,10,5,34,17,-7,-2,-10,9,5,-2,4,-3,2,28,28,-3,-5,-9,8,-6,-5,-83,-14,-6,-22,-19,-33,0,8,-16,14,-35,-2,-36,14,3,35,28,-10,6,2,8,27,7,-19,-7,-30,-9,0,36,21,-22,3,-8,5,-105,-12,28,2,20,-6,15,-4,55,-10,-1,-11,56,35,30,-11,-14,-8,13,9,-34,-8,5,3,6},
{24,-80,0,8,-12,1,-3,32,-5,10,2,-92,-6,-22,28,41,-1,12,12,-7,-6,13,11,-33,-50,5,6,7,-68,2,4,-1,46,56,-11,-52,22,3,17,-21,20,4,-16,7,-1,51,-11,10,-4,15,-23,-36,18,5,1,-14,-3,2,-27,-1,-59,47,40,4,-36,9,-63,-2,62,-18,24,-4,-1,-3,-109,53,-26,-18,-9,-10,0,-31,9,29,32,69,27,-1,27,61,-11,-6,3,4,-67,29,12,7,-26,-10,-86,-7,7,16,8,7,36,40,6,11,-16,0,8,13,0,23,29,-12,61,1,-18,11,-3,10,-46,-1,-3,4,15,-5,-12,-35,0,-9,-13,20,-49,-8,-3,7,-1,-48,-54,31,-1,26,12,-9,27,-5,-9,13,2,-47,12,-6,44,-42,8,-21,38,2,22,4,1,-6,0,-4,100,20,-21,-22,12,0,0,-37,-15,10,10,24,-14,9,0,15,-1,13,-34,20,27,45,-74,11,-11,0,0,-2,35,-5,-3,-59},
{42,3,-6,11,11,15,3,17,-1,-23,2,-19,57,27,-1,11,-8,-32,5,1,-2,7,8,-8,1,15,-17,6,-24,49,0,11,65,34,-10,7,16,-13,-13,-18,13,1,-41,0,-10,-6,2,4,4,-8,3,-37,-51,28,0,7,-33,-1,-42,-23,-29,-34,-42,-13,14,-32,-48,-27,56,-6,13,-24,7,13,-28,4,-12,-41,-5,-10,4,-19,29,-27,41,12,59,4,47,28,6,30,24,0,-5,29,-3,31,-10,22,-16,-4,-39,16,-6,0,-4,33,-10,-35,-23,4,8,32,-7,28,18,-77,40,-49,-21,0,16,-6,-15,-5,-33,-2,-16,-5,-3,-45,7,-63,-5,22,-43,3,2,8,4,4,-27,11,40,24,5,-1,25,-13,-27,4,0,-27,-3,6,48,-28,16,-38,-3,4,15,3,14,-7,-6,-11,96,-22,-42,-8,16,0,1,41,15,-10,5,-19,-8,1,-1,-75,11,19,47,52,11,27,10,22,-3,-22,3,5,44,0,9,-133},
{-7,17,7,9,-37,-5,-13,-1,-20,-11,-1,-4,46,51,-47,7,-2,-42,14,0,-8,2,-3,-23,35,7,-2,8,11,38,-4,15,14,10,-10,32,-15,-13,-7,-13,-3,5,10,-9,-25,-20,-37,-4,1,-30,-17,-55,-50,-7,-5,36,-60,4,-7,-41,40,21,-46,-5,24,-35,-37,-38,23,3,0,-44,9,-6,-4,20,7,-34,8,-5,-5,5,-15,0,26,-13,-13,-10,54,48,22,3,23,-1,-9,-7,-9,18,-1,-6,25,13,-57,17,4,9,-16,70,1,-12,-17,-7,-5,-13,-7,4,8,27,7,-62,-18,-5,36,-7,5,-5,-63,-28,-19,-2,0,-14,7,-43,-7,51,14,-9,5,-5,-3,-24,11,-7,19,8,2,7,8,13,-8,-2,-5,3,-13,6,44,0,7,-19,32,6,31,4,2,-4,-16,29,77,6,-3,21,12,0,2,58,7,5,-7,-11,-23,0,2,-18,18,26,12,67,-8,28,47,34,-7,-67,-10,-15,3,28,7,-38},
{-18,17,2,10,-23,2,-4,-20,-22,-42,-1,-11,0,24,3,25,-6,-18,47,-5,2,-14,3,-26,40,-11,-4,-1,17,1,7,-13,-50,0,-27,0,26,0,4,-25,-24,-6,35,3,-26,0,-21,0,2,-27,-39,-26,13,-26,31,55,-39,-4,15,-16,81,30,-13,10,15,14,-2,-12,-10,16,-1,-34,-3,-14,4,5,7,1,33,14,6,-27,13,27,13,7,-12,3,33,-6,15,10,-13,3,22,-23,2,29,0,-14,33,23,-16,-13,-7,-3,-11,-9,9,0,-2,-6,-1,-73,2,-8,-46,90,0,-19,-20,10,25,2,0,0,-38,14,-17,-5,-2,-11,7,-18,-19,-2,52,1,-2,7,3,31,17,30,-34,1,15,4,-23,-15,-18,-33,-6,27,13,4,-45,1,-3,3,29,-4,16,-5,22,0,-6,99,11,-17,3,13,9,0,8,5,-18,17,0,7,15,0,-6,22,9,5,-62,6,-15,25,18,21,-2,-33,-3,-6,-7,6,10,36},
{-21,0,-3,-10,24,-25,-14,7,44,-40,-9,9,-15,5,27,-41,11,24,21,1,8,2,-6,30,-15,-8,-24,5,42,-25,2,-73,-54,-29,-9,-2,33,1,-63,-17,-37,-3,36,-3,-9,-14,-2,6,7,2,-17,35,43,16,20,11,-15,0,-27,1,98,-27,-9,4,0,41,0,-2,-15,-14,-13,-21,22,-14,6,-16,-29,-30,-6,21,5,-48,-17,1,9,-19,39,8,-26,-7,6,-11,10,11,30,-10,5,-17,20,36,12,0,28,-53,5,8,-2,-73,21,-41,-16,-11,33,-57,7,23,16,32,-19,-5,1,-10,-40,16,24,2,39,32,-15,8,-4,-20,4,-49,11,-53,88,-11,5,-2,7,74,35,25,-51,-26,15,-2,2,-6,-34,-6,5,-18,2,-3,11,15,3,35,9,4,-19,2,12,2,15,15,-6,-58,-23,4,-2,-7,3,-22,-11,11,-5,10,46,8,1,41,-21,27,-54,7,27,-22,-13,-12,-3,67,-2,-17,10,-34,-3,49},
{3,-23,2,-18,27,-33,-2,12,56,-22,7,11,4,0,23,-50,3,-13,-48,-4,-5,-1,-2,48,-64,7,-27,-4,73,-41,-8,-16,-38,3,11,-17,19,19,-63,-18,27,-4,52,-3,-14,-21,-40,4,-3,-36,-18,-27,50,16,-1,-55,-25,1,22,12,-14,-83,21,-9,-28,27,-9,25,-13,-11,-10,1,-57,-4,-11,-24,-53,-2,-35,-13,7,-31,-46,20,6,-21,1,7,-46,14,-11,-48,45,1,0,-21,5,-73,58,40,-15,-10,14,19,-1,1,2,-14,4,-31,0,8,5,18,3,33,65,-1,-29,-5,0,-5,-13,41,-21,-5,42,14,-2,-1,-8,5,-6,-40,16,-79,40,-4,0,-1,7,65,21,-17,-61,-18,-42,10,24,0,-29,-22,-6,-39,-66,6,93,14,-12,30,24,0,-30,-2,4,-5,31,-30,-37,-52,-52,9,-47,0,0,16,18,-2,4,8,49,17,2,47,-19,-31,0,8,37,-40,22,-5,-8,54,-13,-43,35,-2,2,13},
{7,-1,0,-14,7,20,-9,-4,11,-19,2,49,9,-4,15,-42,0,-17,-50,-8,7,-5,0,52,-72,12,-23,-1,41,-56,-6,9,-15,-33,3,-34,-24,1,-35,15,-5,1,44,-4,-34,-19,-73,4,-1,-32,-14,-115,35,-18,-7,-47,-52,7,-1,-9,-78,-92,-8,-11,-17,2,-21,19,-10,-8,-24,-2,-43,-5,-10,-45,-110,-15,-37,-18,2,0,-7,31,0,-15,-6,0,-31,29,-44,-89,50,-6,-39,58,-6,-32,39,1,12,-21,-16,42,3,2,-6,38,-4,9,21,4,-28,61,6,32,81,29,-12,-12,-2,1,22,46,-6,8,15,-11,-10,0,0,12,1,-16,-14,4,18,0,-6,3,8,10,21,-69,-25,-46,-14,5,30,-20,-19,-55,6,-13,-47,-2,82,12,-7,8,-10,5,-28,-8,-19,5,-4,-60,-39,10,-23,-11,-9,-8,5,26,16,5,-8,-16,27,14,-3,32,-17,-35,20,45,16,-24,49,12,-3,53,0,-46,43,-13,0,10},
{18,-23,-2,-13,20,35,5,-7,-42,-26,0,15,5,-53,16,20,-2,-33,-16,6,-2,4,-12,5,-57,12,-4,-9,-3,-15,3,25,6,-26,-17,-14,-27,-12,-15,29,-20,-5,8,-6,-26,-17,-44,-4,1,10,16,-83,3,-6,-2,-15,-91,-9,-19,-4,-55,-79,0,-9,-6,-23,-9,2,-2,0,-12,7,-19,1,-61,23,-300,-47,-24,-17,4,-15,14,6,9,-7,3,-3,-17,3,-5,-42,22,-8,-11,13,-8,5,1,-45,22,-22,-6,46,-7,4,-9,60,-6,29,27,1,-15,37,3,32,51,66,-15,-13,-22,-4,8,6,22,0,14,-22,-36,0,0,16,-4,-17,-23,73,15,-2,-3,0,8,-17,2,-27,-20,-65,4,-14,3,-40,-8,-64,4,-33,3,0,16,7,0,-4,-46,-1,-16,5,-20,1,-53,-7,-9,41,-9,-18,27,-7,2,41,20,-30,-4,-16,5,-22,-2,9,-38,7,-19,59,-11,-2,29,-10,-1,20,-4,0,20,20,-4,4},
{-11,-45,6,-27,11,-2,1,-11,-18,-65,6,16,-29,-55,-6,21,-28,-15,-2,6,-10,4,-4,-19,-51,-3,-14,-8,-12,-11,2,54,-1,-6,-10,-9,-17,-14,-16,-1,-26,-4,-22,-18,-9,-11,15,6,-1,-6,-1,-27,9,-1,-11,-26,-32,-9,-3,-5,-25,55,39,-4,0,-26,-25,0,-2,-2,-6,-10,15,-9,-29,7,-141,-56,13,10,3,-44,-20,0,-61,-30,-3,-6,-29,-28,-6,-100,3,-12,-39,-57,-19,14,4,-41,1,-19,-12,18,2,-2,-6,27,-70,17,16,1,0,17,-7,-1,40,50,14,-37,-4,-8,-26,9,5,-5,3,-18,-8,-3,5,11,-8,49,-2,56,-17,0,-7,4,-8,-66,18,-7,-17,3,-10,-12,-25,4,13,-19,-6,-8,-9,-4,33,10,34,-34,-39,-7,-16,1,-13,5,24,-27,8,58,0,-3,29,-1,-4,21,2,-42,3,-28,37,-85,3,15,-57,-5,-16,48,-2,-6,8,-20,-26,-16,-9,7,-8,9,-7,1},
{-8,8,7,-12,-22,-39,0,-22,-6,-7,0,28,-11,-19,-192,-37,-4,-16,-80,-5,7,0,-4,8,-18,-10,-4,1,38,-31,-1,11,9,-27,5,-17,-6,-107,-34,4,-58,-8,1,4,-4,9,-21,7,-5,-15,-26,3,-46,-2,-7,-28,-12,-2,-27,-9,-41,48,-40,-13,0,-19,-1,1,4,-32,-11,1,-20,3,-20,-21,2,-59,-11,-7,4,3,-23,-21,-191,-8,0,-5,-7,7,-38,-528,-33,0,2,-12,-19,5,-4,0,10,2,4,-7,-1,6,-13,-41,19,-6,-15,-9,0,-8,-12,-6,-11,-5,-18,-11,-11,-7,1,4,-19,4,1,-40,-15,1,-4,-88,-5,-5,2,-9,-13,-3,-7,-7,0,-1,-1,-28,10,-13,-20,-7,-6,0,8,18,-8,-62,-71,-4,31,-18,2,-21,-92,-1,2,4,-27,6,19,-41,0,0,-2,-21,-3,8,0,-10,1,-16,6,-15,0,-15,-3,-32,-33,-12,1,56,7,3,12,12,-13,21,-3,-53,-5,-11,3,26},
{0,-11,4,-14,-12,-13,-14,-45,8,-1,-10,42,1,15,-39,-66,-6,-10,-73,2,-9,5,0,21,-17,2,-8,0,24,-37,0,1,14,1,35,-52,-42,-54,-31,-15,-46,0,-6,2,10,-4,-20,0,-6,-14,-31,-14,-34,18,-15,-24,-7,-8,-10,-6,-9,-106,-55,-44,-3,-4,-44,3,-4,-36,0,-5,-17,3,-40,-7,10,-28,-22,-22,-3,-5,-10,19,-66,-54,36,1,-24,4,-35,3,8,-7,11,-4,-20,-42,6,-1,37,-8,-17,0,-2,-11,-12,-16,11,-3,17,-7,1,33,3,8,45,5,-3,-14,-11,-10,-10,6,-31,6,-7,-16,8,3,8,0,6,-74,44,0,38,3,0,-7,0,19,12,-22,-16,-3,4,-7,29,-1,-24,-57,-2,-38,-47,-15,43,-3,-2,-2,-31,5,-1,-3,10,-7,-63,-42,30,-4,-3,-14,-13,-2,1,-1,-8,-28,-1,-23,9,-7,-5,22,-14,-8,-6,32,1,8,20,-16,-2,19,0,-49,-1,0,-3,25},
{7,12,7,-5,14,8,-29,-47,24,0,3,114,9,20,-7,-90,-11,-5,-47,-8,-2,-5,13,25,-9,-2,-6,8,41,-51,5,15,57,-52,37,-22,-84,-26,-48,29,-24,7,-13,-2,2,-3,-10,0,2,-10,-13,-89,-14,-14,0,0,-29,4,-19,-10,12,-196,-45,-99,-17,19,-26,26,9,-16,-9,19,-3,13,-68,-26,-25,20,-36,-3,0,-22,11,17,-5,8,7,2,-35,14,-23,-70,-3,-14,10,-14,2,-61,-22,15,29,4,10,-7,-2,-8,-11,4,12,1,36,11,10,59,-6,-4,86,12,18,-2,20,-8,22,14,-42,3,28,0,4,-1,-2,0,-8,-19,23,0,36,-5,-8,7,4,12,-20,-54,-29,-59,33,-11,32,15,-31,-63,-8,-12,-52,-2,29,38,9,2,-45,-1,25,-4,-27,-7,-59,-40,19,30,-53,-3,-5,2,1,-25,8,-25,8,-33,16,18,6,70,-13,-26,-32,56,13,-3,44,12,-9,14,-4,-77,-3,5,-3,10},
{0,-14,5,-5,5,25,-5,-24,11,-19,0,63,29,-7,0,-33,9,28,-16,1,-6,5,8,18,-50,-4,-30,12,-18,-147,5,-14,14,-45,-1,-9,-44,-20,-20,11,-9,4,32,-2,-50,7,-8,6,0,-3,-20,-144,19,-11,2,-2,-5,4,8,4,17,-47,-18,-67,-12,28,-42,16,41,10,17,6,1,-9,-77,7,-51,31,-53,-1,7,-39,-18,77,3,115,-27,-4,-23,41,-39,-80,3,-2,2,-12,0,-31,-22,7,19,-12,15,-4,-6,7,1,21,33,4,44,11,-9,43,-11,-6,84,57,28,14,0,5,40,16,-13,1,26,4,9,8,-2,-13,0,6,30,6,22,6,3,-9,1,-34,-17,-27,-28,-23,-10,-2,32,9,-30,-64,6,-9,-27,-5,33,49,0,20,-33,2,10,7,-26,-5,-96,-24,-29,-21,-13,-19,7,4,-8,-39,0,31,7,2,-20,5,-11,54,-15,3,-10,64,23,3,-1,-24,-8,1,0,-70,-11,1,4,13},
{19,-61,6,-8,-1,8,0,-28,-5,18,5,-42,-21,-21,7,24,-6,38,46,6,7,2,5,-22,-96,-15,24,-4,-45,-92,-2,-10,2,8,7,-12,-15,-1,44,-11,19,-3,-5,4,-32,46,-9,-3,-5,-11,-27,-55,11,-37,24,-42,-9,0,14,28,-16,73,52,-28,-22,7,-60,-2,62,-3,34,-5,14,-5,-133,46,-32,32,1,0,-7,-53,-23,132,34,114,-7,-3,13,78,-37,-53,22,10,-44,28,-11,-24,-4,-37,-29,-18,25,13,6,-8,40,41,17,16,17,1,-5,27,-7,1,25,6,65,0,-2,-3,8,33,-1,-1,11,-8,20,-4,-1,-52,10,47,11,1,-44,0,0,-7,-2,-19,-26,21,-11,13,-11,3,16,-17,0,29,-4,-7,27,0,16,0,-1,-12,4,-6,36,5,4,2,-55,12,37,12,-3,-27,-2,0,8,-118,-27,24,-2,33,-22,20,2,8,3,23,-27,64,16,14,-63,-15,0,-30,14,-66,-4,8,-2,-11},
{41,-30,-3,3,-23,0,-2,-5,6,9,-2,-74,27,0,-2,51,0,3,21,-4,5,-6,6,-27,-27,1,20,1,-63,-29,2,22,39,53,19,-29,14,4,37,-55,22,-7,-24,7,-25,47,-8,5,8,-10,-28,-44,-27,0,-7,-35,-30,-3,5,-23,-18,49,56,28,-5,-1,-69,-11,88,-18,27,-19,18,0,-107,39,-33,-10,32,-9,-1,-18,20,-15,59,67,14,-9,37,95,14,-9,26,-5,-24,-13,-3,33,-11,-2,-38,-18,0,7,7,6,-1,-5,-2,11,-38,0,-9,14,-3,1,-19,-54,44,-15,-8,2,-42,22,-34,0,-24,-20,8,-2,0,-47,-1,1,0,19,-62,-1,3,-4,-2,3,-45,16,11,25,17,2,24,-3,-9,16,-3,-10,27,2,0,-39,0,3,57,-1,39,-4,35,6,-12,-7,113,36,-10,3,22,-7,-1,16,-38,14,8,2,8,11,5,-52,28,-1,-7,43,16,23,-75,-24,4,-40,6,-27,41,6,-4,-68},
{12,14,-2,-26,-10,0,1,-8,-23,38,11,-41,42,25,-23,-1,0,-51,38,-2,-2,0,9,-17,18,11,17,5,-13,24,5,42,58,12,-8,-5,31,19,23,-24,-5,-6,-13,0,-21,-27,-22,-5,2,-12,-24,-15,-68,20,-19,20,-40,0,20,-34,16,-10,-13,11,37,-16,-45,-2,49,-6,7,-21,2,1,-64,2,0,4,18,-2,1,0,37,-4,50,-22,-25,11,32,72,4,3,47,3,53,-11,-7,34,-23,1,-6,-26,-36,12,-7,0,4,31,-12,-9,-46,-2,14,6,0,-2,-41,-35,1,-25,-25,-6,-4,4,13,-6,-42,0,-28,4,-5,-12,0,-23,-1,32,-11,-12,0,3,-8,22,-11,8,47,-3,5,-16,9,22,-5,3,4,2,10,6,-29,4,4,-36,52,-6,11,-6,38,-5,-29,6,60,0,-14,13,23,-6,7,35,-16,43,-2,-28,0,10,13,-73,17,-3,69,56,-6,5,3,-1,5,-47,7,-11,21,11,8,-75},
{-14,29,1,-12,-4,14,-3,-37,-25,53,4,-3,3,33,-12,2,-6,-33,32,6,1,-4,-12,-38,40,-3,33,4,-4,-5,4,35,6,4,-20,-7,5,19,61,-11,-30,-4,19,0,-18,-3,-26,3,-4,-4,-43,-22,-54,-24,-17,26,-51,4,49,-34,11,8,25,31,1,6,-16,0,10,-4,-8,-24,-20,1,-40,8,0,52,45,-23,-6,-2,45,70,32,-8,-46,3,30,52,0,29,30,-1,15,-4,-2,50,-12,-13,3,-6,-26,1,9,-1,11,1,-3,6,-5,-4,-8,-34,6,-1,-93,37,0,-10,-32,-10,11,6,29,-6,-46,1,-18,-6,-1,0,0,7,-8,57,15,-5,-2,-2,1,30,13,24,21,-35,4,8,-12,-8,6,2,-3,15,28,-5,-63,-8,7,-20,50,2,27,0,25,-3,-28,58,12,7,15,6,22,2,0,18,-8,45,0,0,-11,0,2,5,34,-8,-7,2,-8,4,-5,-13,0,-54,-14,-16,5,14,1,-4},
{-27,4,-7,-1,24,36,-8,-9,-7,28,-12,32,-56,19,13,-7,1,-2,30,-2,-1,-12,-6,-42,27,-28,3,8,-9,-6,1,0,-36,-10,-4,-4,13,16,71,-6,-49,0,12,7,1,5,13,2,0,25,-14,8,-15,-38,7,18,-29,2,14,-24,17,-61,6,29,14,26,22,-20,-35,8,8,-26,17,3,8,22,-39,21,46,1,5,-24,26,42,61,4,4,-1,12,43,2,45,41,-11,-10,36,-10,28,-21,0,7,-22,-3,-35,6,-7,10,-9,7,-21,46,0,-9,-71,4,19,-79,49,-35,6,-3,13,-22,23,25,5,0,5,-25,1,-3,-27,7,-15,-18,29,46,-4,-1,0,6,61,13,17,-18,-32,6,-5,-36,-28,19,-14,8,15,31,-11,-88,-16,0,9,29,0,-11,0,28,6,-29,64,-10,-33,-21,30,7,7,1,-23,-13,51,-3,33,-9,5,-6,20,59,-14,-62,38,3,-1,-23,-13,-9,-21,0,11,-1,3,3,9},
{-15,-13,6,16,20,9,-1,-2,49,36,-4,32,-18,0,18,-92,7,22,-4,1,1,1,-7,16,-50,-28,-2,-2,15,-50,-6,-38,-24,-6,36,25,26,4,-19,-15,-57,4,7,2,-31,-18,2,5,0,25,-19,18,0,20,13,-53,0,-6,-7,27,58,-87,-31,8,2,29,-4,-4,-12,-11,8,-14,30,-7,-19,33,-77,-45,19,-15,-5,-36,-3,-4,27,42,59,3,-32,33,-40,-8,77,4,44,-11,10,-41,15,35,-8,-10,9,-33,-1,0,0,-17,10,-66,15,-3,30,-18,2,55,39,12,-74,9,0,10,-44,15,20,2,47,9,-25,-1,2,-43,10,-19,15,12,41,4,5,5,3,42,35,-7,-50,-18,0,8,10,-9,-19,-17,5,-22,-8,-3,41,-20,-12,44,7,-8,1,2,9,-2,-3,-50,32,-33,-30,16,-18,1,-8,-36,29,29,8,7,40,13,-5,28,17,-5,-36,32,34,-26,21,-25,-5,48,1,-18,0,1,8,13},
{-3,-23,0,-42,3,-35,5,-5,96,27,-3,22,-8,6,18,-69,-2,6,-13,-6,-6,3,4,32,-97,-5,-25,8,-8,-81,0,-24,-13,53,33,6,8,10,4,-17,4,2,26,0,-11,21,-27,-3,8,-28,-16,-27,2,-6,-8,-112,-35,3,30,32,-40,-36,29,-16,-49,9,-22,9,26,-29,5,-2,-48,6,-42,0,-57,-4,19,-45,0,-25,-26,23,13,93,25,8,-9,45,-53,-56,71,2,14,0,2,-83,40,10,-20,-12,0,39,-5,-2,11,15,-5,-17,11,8,1,27,5,44,91,-1,-47,4,-8,-9,-40,18,-16,-9,27,-19,6,3,-6,-10,5,-12,23,-27,1,7,-7,-6,-6,36,19,-6,-76,-10,-55,6,36,-2,7,-1,-4,-17,-14,4,98,-34,-19,12,23,-7,0,6,-2,-6,24,-46,10,-36,-21,20,-61,4,0,-28,39,0,0,-12,51,9,10,7,5,-20,0,12,45,-19,21,-24,-3,21,14,-71,16,9,0,-11},
{-3,-5,7,-42,17,17,-9,-15,-3,0,-2,47,4,4,13,-49,-3,-20,-41,-1,0,-3,-1,28,-88,-1,-47,7,-23,-114,5,-17,3,-6,-10,-20,-33,0,-11,12,46,0,24,2,-13,26,-21,5,-6,-30,5,-147,12,-29,-12,-50,-61,6,0,-4,-63,-36,11,-6,-41,10,-14,31,20,-21,-18,-6,-57,3,-8,-37,-76,4,33,-29,-6,-24,-11,47,22,69,0,0,7,52,-46,-64,67,-2,-19,66,-17,-15,-1,1,18,-36,-17,45,6,1,12,50,0,27,37,15,-15,72,-9,23,62,24,-11,5,-9,-14,18,18,-20,9,15,-9,-11,2,0,21,-2,0,-36,4,-12,10,-1,-2,4,-6,15,-32,-17,-19,-28,-1,22,0,-9,-50,-3,7,-32,-3,58,-11,8,-4,2,-5,-30,3,-23,5,-37,-6,-42,-20,-1,5,-7,-7,6,15,18,-14,2,8,20,-1,11,8,2,-27,-11,27,-1,-11,23,-1,-2,41,10,-63,27,5,-2,-1},
{-7,25,-1,-19,29,26,-14,-5,-55,-41,-3,37,-5,-20,-9,-2,0,-57,-7,8,-2,9,-5,8,-50,8,-15,1,-37,-28,-5,17,18,-36,-26,-20,-33,-13,-8,40,35,7,16,-5,0,-4,-5,-8,-3,-16,15,-149,-7,-19,-14,21,-75,-1,-30,-16,-91,-25,1,14,-34,0,-8,18,-10,9,-14,-6,-19,-9,-29,-9,-158,-54,12,-6,3,-39,25,8,3,40,-15,0,-24,16,-3,-69,55,-10,-74,22,-12,31,-22,-45,28,-14,-15,-43,-8,0,15,27,7,29,66,-6,-20,44,-8,3,22,35,-2,-1,-7,-8,19,8,2,0,21,9,-33,0,-11,21,-4,0,-65,30,0,-4,5,-5,3,-31,-14,-9,0,-40,25,11,1,-33,-15,-44,5,-8,10,-7,15,7,5,-5,-32,0,-65,-5,-43,8,-96,19,-13,1,0,-8,21,-9,0,6,21,-30,3,20,7,10,1,-12,-6,2,-56,41,-55,-9,17,-1,-4,19,-5,-6,34,10,-4,-3},
{-44,-28,5,-3,28,1,-40,3,6,-51,-5,10,-21,-42,-18,17,-10,-17,17,8,-7,0,-5,-15,-51,-2,-30,-9,-46,11,7,62,-6,5,-25,-18,-11,-21,-2,18,-11,6,-17,-42,4,-31,2,-7,-3,-11,4,-44,-56,9,-10,-24,-26,-10,-25,-5,-37,62,29,-20,-41,-44,-5,-20,-9,0,-11,-25,10,-1,57,22,-90,-41,13,-14,-4,-65,-14,-60,-67,-21,13,-12,-19,-22,7,-54,8,1,-48,-15,-21,12,0,-72,-2,-36,-23,-27,-1,1,-9,-1,-25,23,20,-16,-20,28,-12,-5,20,-7,-11,-48,11,5,-17,12,1,3,19,7,-8,-1,4,23,-4,16,-18,27,-22,-11,-4,-8,-8,-44,2,22,4,25,-2,0,-16,-24,18,1,3,-8,7,-8,35,2,9,-49,-6,-3,-35,-4,-37,8,25,-12,19,12,-4,8,18,-8,5,30,3,-31,0,-21,27,-41,6,5,-21,18,-68,63,-31,7,9,-17,-15,-12,0,31,-8,-10,2,-1},
{-12,3,0,-31,0,-11,0,21,-1,-3,-6,29,-12,-7,-61,-103,-18,-41,5,-5,0,0,3,-16,-31,1,-14,-4,-3,-97,1,-28,-74,-6,10,1,14,-48,-1,11,-45,2,-14,-9,19,-42,-59,6,-3,9,-27,-40,-56,0,-45,-30,-30,-4,-37,-2,-10,29,-47,1,-13,0,26,14,-11,-115,-29,20,-20,0,40,3,9,-56,-368,-15,5,-33,8,-164,-288,-35,-14,5,-35,0,-69,-51,3,-8,-1,2,-8,7,48,10,-717,-2,13,-6,-7,3,-32,-17,0,7,-26,-15,0,-25,2,-55,-374,9,13,-18,11,-15,7,34,-13,0,-26,7,7,1,7,-60,-6,33,6,-2,-38,-4,-2,-3,4,-38,-18,14,16,17,-4,-20,-162,1,-1,27,6,-34,-17,-2,-28,22,5,-10,2,-4,-13,-7,-1,8,-12,-45,5,0,2,-28,-3,3,-8,-39,-21,-10,-6,-70,5,29,0,17,-12,-1,-6,-17,-1,-65,16,19,-27,-27,-5,-12,-2,-9,-1,-292},
{6,18,-8,-27,-13,-20,-29,13,9,15,-2,29,18,0,-4,-108,7,-27,-16,2,-3,-11,-8,25,-34,4,4,-6,42,-50,1,3,-22,-12,-6,-31,-2,-45,-27,2,-78,6,-10,-2,17,-13,-50,5,-10,-39,-59,-73,-22,-20,-28,-15,-38,-1,3,-22,-2,-8,-29,-29,-17,-9,-43,45,-3,-43,-5,-18,-36,-6,-10,-51,3,-9,-11,-12,7,-18,11,3,-74,-72,33,-8,-35,32,-64,34,27,-5,17,4,-20,-24,25,4,24,7,-2,-3,7,-12,0,-12,10,9,-30,-1,2,45,5,7,-23,6,1,-25,-13,-24,10,27,-51,7,34,-4,5,-2,-9,-23,5,-89,11,-13,32,4,5,-7,8,-1,-18,1,6,-4,-12,-4,18,-8,-74,13,-9,-42,-33,-11,51,-5,-8,-22,18,-5,-31,-4,-27,0,27,-44,11,30,-50,-26,-39,3,0,-11,-13,-5,-4,-24,5,43,-2,17,-19,-45,9,1,4,10,56,4,-6,20,0,-72,6,-24,-3,36},
{11,24,2,-16,-5,17,-3,-4,-2,1,-5,61,23,14,23,-97,-4,-14,-33,1,-7,-5,-6,45,-48,-8,-25,-1,42,-56,-5,11,14,-33,1,-21,-21,-23,-45,29,-6,-3,-6,-8,20,-59,-13,-1,6,-46,-23,-128,7,-9,-18,2,-9,-2,-19,-16,-5,-180,-22,-49,-26,4,-31,58,15,-12,-16,6,-8,1,-42,-44,-47,5,-78,0,-8,-23,21,14,-16,23,17,1,-52,36,-19,18,45,9,9,19,-5,-20,-1,5,24,5,3,-15,3,-4,5,-14,25,29,20,15,3,78,9,-4,37,26,13,-12,22,1,22,13,-50,7,50,-5,-4,-9,-11,-9,6,-15,9,3,28,-4,-4,-3,-6,-1,-22,-58,27,-57,15,-5,22,7,-25,-26,5,-19,-49,-6,30,29,-12,-20,-16,-2,-45,-5,-35,7,-108,-51,10,38,-59,-15,-15,3,5,-11,0,-23,-1,-17,0,24,4,21,-15,-32,-8,43,14,9,17,-3,-2,30,0,-80,19,-8,4,21},
{-8,6,-8,-26,3,5,-5,-11,-1,0,-5,38,9,9,31,-54,13,24,-28,1,2,-10,-3,23,-91,-10,-22,10,-14,-89,-1,-16,1,-29,15,10,-9,-4,-20,7,23,5,3,-10,-1,-1,7,-1,4,-29,-17,-140,21,-41,0,0,11,-1,-2,16,0,-64,-5,-42,-17,13,-18,4,31,-5,5,12,2,0,-75,-10,-57,16,-88,3,8,-72,-19,58,-33,124,-4,-12,-34,47,-32,5,42,1,10,17,1,-37,-5,-8,24,-11,12,-10,-2,-5,0,1,40,21,39,0,-4,62,0,-4,26,24,0,10,17,-13,11,3,-12,7,48,4,2,0,-4,-5,3,26,18,8,37,-3,-6,-3,-8,-27,-16,-35,8,-16,7,-1,34,1,-13,5,-10,0,-41,0,27,30,1,5,-22,3,-37,-8,-18,6,-118,-16,-26,-46,-30,-15,-6,7,-4,-24,16,3,-1,14,-23,0,10,28,-23,-20,-35,48,19,0,-25,-9,0,15,0,-78,0,10,7,38},
{-3,-19,-5,-2,-27,-26,9,-14,-23,-20,-2,-34,-37,1,36,16,-4,39,28,-5,-1,-10,4,-8,-84,2,-2,3,-42,-64,8,-12,0,44,14,24,-7,7,19,-17,29,1,-9,-8,0,44,5,-1,1,-3,-22,-13,13,-8,11,-60,12,5,-3,36,27,46,67,0,3,5,-20,-32,47,-4,19,-1,26,-11,-95,40,-38,6,-20,0,0,-96,-34,57,1,104,45,2,1,51,-16,17,42,11,-19,-6,-6,-12,22,-32,-22,-3,20,45,2,-1,25,-18,23,13,-6,-7,-29,-1,8,-19,-25,2,38,-4,13,0,-44,23,11,-2,9,-6,19,4,-3,-43,5,47,15,-13,-6,1,1,4,4,18,-8,5,2,38,-7,4,21,-2,7,33,3,33,-4,12,15,7,-16,1,2,0,9,4,30,1,-44,30,28,-12,-4,-17,-32,1,5,-41,-7,-6,0,25,-32,-28,-5,-16,-7,-12,-68,19,34,-13,-75,-13,0,-40,-9,-66,-20,14,3,-18},
{22,8,-2,26,-34,-4,-6,-22,-24,-25,4,-58,24,10,22,37,0,-8,30,-2,0,-10,2,-19,12,23,33,0,-38,-40,5,45,22,21,22,1,13,40,14,-21,7,-7,-9,-8,-5,-17,-24,3,0,10,-12,14,-14,11,-9,-23,5,-7,-6,-7,66,10,68,32,18,-9,-20,-23,34,-2,18,-7,39,-10,-57,25,-47,-21,5,-2,-2,0,12,-73,-1,26,9,0,-11,33,60,3,19,-4,56,-56,-2,21,19,-9,0,0,-21,60,2,-3,-6,-19,0,-14,-42,-2,-28,-49,0,-19,-37,-43,-15,-10,-18,-4,-74,38,23,-5,-36,-22,1,-1,-3,-29,0,32,8,-10,-43,0,-6,2,-1,43,4,-2,19,18,43,-5,10,23,9,18,-2,48,7,4,-25,18,-14,21,39,1,11,-1,46,-4,-5,-11,15,22,9,19,-3,2,0,72,5,1,-2,-14,-19,-27,5,-69,-10,8,-15,44,1,-21,-63,-27,-9,-58,-1,-1,-3,24,-3,-39},
{-16,48,-5,-7,-14,13,-8,-26,-38,-1,-4,-36,21,15,16,26,-1,-40,16,1,-3,3,-5,-9,18,27,40,-5,-2,-1,0,55,50,-6,-14,-38,15,23,23,-1,-12,-6,9,-4,1,-17,-34,-1,-9,32,-9,7,14,15,-18,25,-6,-8,20,-48,39,1,80,21,2,-12,-22,16,11,-3,20,14,-8,-8,-38,-9,-21,37,7,5,2,11,28,12,-40,-37,-49,5,-28,16,24,-24,10,11,56,-16,-9,48,3,-18,30,-7,-20,17,0,2,15,-26,-8,4,-39,-6,-7,-34,7,-16,-44,7,1,-16,-29,-22,21,11,32,7,-36,-2,4,5,4,13,-3,18,3,11,-17,0,7,-6,0,51,-5,4,41,-17,24,16,-18,4,-2,14,-7,47,7,5,-55,45,9,-24,20,0,-6,-5,30,1,-32,14,-1,1,24,25,24,0,4,38,13,26,-2,0,-43,-24,5,-52,-20,-7,18,17,0,-41,-55,-11,-12,-70,-4,26,-12,-2,-6,-54},
{-32,43,-5,-7,-13,23,0,-14,-24,13,-10,15,-55,9,19,39,-3,-8,-2,1,3,4,1,2,6,32,7,2,-4,7,1,31,18,6,-22,-50,-14,20,52,1,-19,8,8,10,8,10,0,7,-2,25,-5,28,22,16,-8,2,0,-4,20,-67,8,14,51,10,-21,0,1,13,-18,4,4,8,-1,-5,18,-12,-17,68,-23,13,5,8,38,66,-11,-43,-17,1,-7,18,-8,12,3,-5,19,39,-6,56,1,-26,27,-12,-10,27,-4,-6,21,-10,-19,31,0,-1,-4,-64,-1,-1,-50,25,36,1,-14,4,1,15,35,-5,-23,-15,13,8,-4,6,-1,22,3,24,5,-6,-3,1,-8,46,-3,-14,16,-40,24,-4,-48,-3,33,-5,5,41,12,6,-72,26,20,-7,17,0,0,-2,21,7,-24,36,-27,-3,24,19,36,-5,-3,14,-2,23,-2,20,-36,-6,1,-1,1,-19,-18,-36,-11,-44,-30,-21,-16,-34,-16,31,-31,2,8,-25},
{-26,26,1,39,-2,28,-6,7,21,50,-3,18,-65,9,10,-6,5,-5,-2,3,6,1,-2,-16,-22,-1,23,2,17,19,7,-5,4,-10,29,-21,-7,17,11,-9,-12,0,-13,18,-8,-12,30,-7,4,33,7,10,-7,4,4,-5,17,-4,18,-34,12,-72,19,-1,12,18,5,-2,-40,47,18,-12,-16,-1,12,16,-25,32,-31,13,-7,-6,16,12,28,-15,-17,2,-23,62,-25,65,28,-11,-3,30,8,20,0,-3,3,-9,-30,-17,-4,0,-13,-10,-3,-32,5,1,5,-52,5,7,-39,-21,2,5,-18,7,-38,25,8,7,-3,-7,-10,0,-4,-19,0,-18,2,23,3,4,-6,-6,-4,17,5,-5,-9,-2,4,-2,-30,-12,-19,-9,-5,22,1,-1,-25,-9,11,24,-3,0,-17,-7,27,3,-1,-3,2,-11,6,18,15,5,1,33,2,36,7,48,-25,13,7,35,30,4,6,42,5,-32,12,-5,-2,0,0,32,-17,10,6,-22},
{21,-3,-4,29,-48,-3,-6,17,44,50,-3,-13,14,0,8,-77,-5,24,-24,5,6,0,-4,26,-63,-28,28,0,0,-57,0,-45,6,24,48,48,20,-7,0,-48,-49,0,-1,1,-27,-22,24,2,9,26,-9,-8,-54,14,0,-76,28,-6,1,2,77,-86,-9,-8,6,21,13,-12,44,-21,46,2,29,11,-29,22,-45,-8,-31,-35,7,-31,2,-58,44,45,71,1,-30,42,-49,14,80,-5,54,14,-3,-36,7,28,-5,0,0,-8,-7,4,-16,-20,-14,-61,-15,0,3,8,-3,39,45,-33,-40,24,-20,14,-51,0,-15,-1,33,2,-2,-2,-3,-56,0,-29,16,57,-4,12,5,-1,-4,22,13,-2,-52,-5,-10,-18,17,10,-22,-12,-3,-2,17,-7,65,-30,-24,19,0,5,18,0,35,-7,48,-90,42,26,-17,4,-32,2,-8,9,-2,27,2,-31,39,15,8,-19,21,-2,-13,-9,25,-10,48,-17,-2,33,-2,-27,12,13,7,-25},
{36,-31,1,-37,-22,-12,0,-8,39,23,-4,-53,-3,6,5,-55,-10,18,6,-2,4,5,-4,30,-79,-24,-5,-2,-50,-102,-5,-23,0,80,52,35,2,0,31,-33,3,-7,0,-14,3,52,-1,5,10,-23,-27,-64,-69,-18,12,-108,-18,-5,16,2,-10,-1,32,-27,-62,0,-3,-6,80,-57,29,-13,-26,-4,-39,11,-14,36,38,-61,8,-58,17,24,10,127,43,-9,21,57,-60,-11,80,-1,11,54,-6,-69,19,2,-15,-27,-11,27,-8,10,30,9,0,-14,29,5,-27,46,-3,44,43,-7,-28,3,-27,8,-50,19,-26,1,36,-22,-12,0,0,4,9,6,23,17,-33,7,-3,0,5,27,9,11,-89,2,-45,-5,45,-1,10,0,-9,-7,12,2,52,-48,-9,-8,18,5,43,-3,22,2,40,-30,48,-29,-18,7,-70,2,6,-39,7,3,-3,-12,40,5,0,-39,10,3,-38,-12,27,10,-5,-21,6,-1,2,-91,14,9,-10,-14},
{-4,10,3,-31,9,18,-11,-23,-8,5,7,15,7,3,1,-8,1,-21,3,7,5,-8,-10,28,-66,-3,-38,4,-84,-122,7,-5,12,9,2,12,-42,-3,0,-6,45,-7,2,-12,9,45,11,-5,3,-48,-13,-133,-27,-38,-6,-25,-32,1,-10,-14,-62,-32,8,11,-69,3,1,23,39,-27,-4,-17,-25,10,20,1,-14,23,41,-44,-5,-70,27,52,21,115,24,0,19,77,-45,-7,63,9,-25,78,-3,7,-32,-26,13,-39,-18,25,-2,-1,44,-2,19,12,77,0,-28,67,-3,21,32,25,-14,3,-8,-9,15,11,-37,6,24,0,-20,-6,4,10,-5,21,-18,20,-15,-6,-1,4,-5,-18,-9,10,-9,11,-26,-1,19,0,-11,-57,4,4,-19,-4,11,-32,10,-16,3,4,-29,0,-8,3,-75,35,-28,-53,-7,-4,-9,-8,-7,17,-2,8,8,22,-2,-12,4,-29,6,-1,-46,5,-8,0,-89,-30,3,8,9,-92,24,23,4,0},
{-6,16,-5,-34,27,19,-26,-9,-62,-49,-4,37,0,14,5,4,6,-46,-19,3,1,4,-2,25,-24,-7,-19,-1,-73,-23,5,24,24,-25,-27,-9,-35,-10,-14,33,60,-4,13,-8,20,-3,-12,-1,6,-39,12,-187,-7,-47,-22,32,-51,-2,-64,-10,-79,-49,-8,9,-75,2,2,39,-13,-4,-14,1,-25,1,-3,-18,-48,-32,13,-1,-1,-64,32,17,0,47,15,-7,-23,16,7,-42,34,-2,-60,22,-8,35,-54,-35,23,-7,-25,10,0,-10,45,15,-1,-5,70,-1,-5,56,-10,-9,-6,52,-5,0,-3,-20,23,5,-19,9,4,13,-38,-6,-4,17,6,-4,-65,17,11,-2,8,-2,-7,2,-18,-2,1,-16,36,-7,5,-17,-20,-54,-5,0,-10,-1,7,4,8,-13,-11,-6,-99,5,-40,-8,-84,25,-18,-36,-9,-11,25,0,5,18,-3,-31,3,39,14,15,-1,-13,-3,-6,-41,34,-74,-15,-15,15,-6,23,-4,-16,33,16,-5,3},
{-35,2,-6,0,10,1,-15,3,-57,-53,-8,-10,18,-19,-31,14,13,-14,6,-8,-3,6,-2,-10,8,4,-43,3,-41,17,0,18,-21,6,-51,9,-26,-10,-3,3,14,8,-11,-64,4,-26,-9,-2,4,-31,-2,-27,-21,2,-8,22,-24,-7,-17,14,-40,46,0,-20,-89,-13,-59,-14,-12,-35,-22,-45,-5,3,23,-3,-39,-22,-14,-60,-4,-78,-4,-37,-98,34,6,6,0,-34,22,27,25,-8,-66,-1,-8,49,-12,-68,-15,-36,-28,-23,5,6,-1,1,-12,-7,-20,-12,-20,9,3,1,-37,-58,27,-27,1,-2,11,13,25,-5,-10,0,-26,-3,3,13,4,14,-25,3,10,3,5,-5,7,6,-8,11,2,0,15,-15,-18,-38,21,-11,-2,-7,-5,0,9,12,-13,-23,3,5,-18,4,-49,7,32,12,5,-51,9,3,42,-4,7,26,13,-6,-1,-27,3,-50,5,-10,3,2,-43,52,-101,-19,5,26,-9,-5,0,22,-15,-53,-4,-19},
{-30,18,-4,-15,-20,-2,-7,0,-5,11,1,-6,2,18,-36,-44,-25,-35,-4,6,-2,-6,-3,-25,-25,-51,-4,6,19,-29,1,-28,-11,-25,-6,-3,16,-62,-100,-10,-42,-8,17,-7,-4,-49,-20,4,1,-36,-22,-23,-23,-10,3,-16,-32,6,-18,5,-9,29,-24,-1,-9,-11,3,21,-15,-9,-41,-48,-36,3,42,-16,12,-25,-13,-13,-1,15,9,-47,-18,-51,-10,-5,-11,24,-58,-717,-20,-11,-49,-35,-27,8,27,8,11,1,-21,-9,7,-9,3,-21,-24,-32,-3,-6,-6,-52,0,-1,-43,3,-18,-39,-2,0,6,9,-11,-10,-40,35,-25,-9,-6,-83,0,-21,-7,9,7,2,-9,-4,-1,25,-2,0,7,-8,-43,-15,-32,25,-28,12,2,-72,-15,0,-14,-31,-17,-63,20,-7,-7,-6,-12,-4,3,-12,-3,9,3,-9,-16,-9,1,-12,-23,13,0,-16,-8,16,0,-12,-39,-7,2,-12,6,4,16,4,-15,1,6,-21,5,-3,-7,12},
{17,23,-8,-42,-11,1,-17,24,2,7,-10,19,22,11,22,-147,-2,-34,1,0,6,4,-6,38,-11,-17,10,-6,31,-69,4,5,-12,-15,-24,6,23,-17,-15,-5,-72,2,22,-4,18,-89,-81,-3,4,-22,-65,-72,-28,-22,-20,-5,-56,4,-10,-36,-21,-48,-16,9,-40,-18,-11,29,-3,-43,-24,-27,-50,1,30,-47,7,20,-8,-32,0,-36,22,2,-62,-69,37,-10,-56,54,-73,102,37,7,4,17,-23,-22,24,-6,19,19,0,-27,0,5,4,-6,1,4,-37,-2,-1,18,-2,35,-99,33,-2,-29,-23,-29,33,16,-52,-2,17,2,-14,4,-3,-30,2,-76,14,7,17,-9,-7,-1,-8,17,-19,-6,-1,-9,-28,-6,15,-3,-87,6,0,-41,-13,-10,45,3,-21,-38,26,-3,-30,-4,0,-1,-2,-36,2,2,-23,-23,-27,-3,3,-25,-36,0,-5,-44,1,48,-4,6,-10,-35,12,-10,26,12,25,15,-16,41,-11,-29,7,-48,6,26},
{4,33,3,-15,-22,18,-7,13,-12,14,4,14,34,0,29,-86,-8,-15,-32,-3,-1,5,0,52,-33,-7,-10,10,8,-36,-6,9,-16,-10,-2,-8,15,-10,-33,19,-12,1,-13,-28,17,-104,-11,-9,0,-25,-47,-115,12,-15,-32,17,10,1,-23,-36,-34,-134,-44,13,-28,-19,-13,38,-15,-20,-36,-14,-20,7,-11,-29,-57,2,-96,-25,6,-68,20,6,-49,10,47,7,-65,51,-5,81,85,2,-5,58,-4,10,-1,-12,44,25,-13,-38,2,-3,3,0,27,41,6,3,-15,79,-6,36,-58,35,-3,-9,4,-9,35,7,-45,0,59,-20,-17,2,-12,-8,-1,4,1,21,50,11,-2,-9,-5,5,-25,-54,32,-35,-1,4,20,0,-42,-18,0,-17,-36,6,39,10,-21,-32,-5,-1,-81,4,-12,-2,-65,-62,32,-13,-36,-26,-20,7,-6,-7,-47,-17,-2,-23,-6,56,4,9,-24,-41,21,16,21,9,23,5,2,40,-6,-47,31,-25,-5,43},
{-4,22,0,-27,2,-16,11,9,-9,-12,-12,0,-10,12,52,-60,-4,-10,-58,0,2,0,1,55,-76,-1,-35,-3,-16,3,6,-30,-4,-14,18,-12,13,0,-33,2,38,1,-15,-24,22,-34,30,1,5,-46,-3,-128,40,-33,-13,31,6,-6,-41,-8,-59,-52,0,2,-12,4,-10,13,0,2,-14,11,-21,0,-50,-12,-48,-25,-61,-15,2,-110,-33,47,-76,50,24,0,-9,50,-31,39,50,7,-21,52,0,-15,3,-13,31,-22,1,-22,6,-1,12,4,48,15,17,8,0,68,6,18,-30,9,5,-2,20,-6,13,4,-64,4,48,-1,-14,-3,-9,14,7,12,5,-10,66,0,1,2,3,-8,-12,-46,10,6,14,-2,30,-4,-5,14,-3,9,-67,-3,43,27,-13,-23,-35,-4,-85,4,12,5,-63,-1,-17,-105,-34,0,-23,-7,5,0,11,-10,3,11,-9,22,-4,-23,-6,-29,-19,22,5,-10,-12,14,18,27,0,-53,22,18,-10,10},
{-34,-7,0,-13,3,-56,15,7,6,6,-1,-29,-51,9,42,-20,3,21,4,-5,-6,-7,4,33,-67,14,6,-12,-49,6,-2,-38,-8,30,14,-15,19,11,-2,-9,24,1,-28,-10,16,18,-3,6,-2,-8,4,11,41,-1,1,-52,9,-5,-23,37,11,1,33,11,-8,-10,23,-55,15,-24,-5,1,15,0,-26,37,-49,-29,2,1,-1,-109,-36,1,-21,61,65,10,19,28,-3,6,23,-3,-10,-9,-7,-9,27,-3,-26,-27,2,43,4,-3,19,-7,13,9,-3,6,-11,8,1,-1,-54,-1,-17,-14,13,-7,-51,20,13,-5,31,-5,-36,6,8,11,-4,10,-11,-23,19,0,2,-2,5,24,-7,6,-3,37,-15,-18,-9,28,19,6,-4,45,-34,4,40,30,-1,-5,-30,-6,-17,-7,27,-5,-29,64,27,-29,-17,17,-25,7,-5,15,54,-37,0,10,24,-39,-7,-33,-8,-7,-69,-31,15,-28,-21,0,0,-4,7,-30,-17,29,3,-12},
{-35,4,3,4,-17,-8,-4,-8,-3,-3,4,-18,-8,-7,32,0,3,-20,26,7,-5,1,0,23,25,41,13,-12,-48,5,6,-6,0,27,13,-36,25,10,-6,-5,-22,6,-28,-13,27,-9,-5,3,0,-13,6,49,43,5,6,-16,1,-1,-15,3,58,-27,62,29,18,-18,17,-22,-2,-8,-5,11,10,0,-2,-3,-64,-31,25,-4,0,12,11,-77,-28,26,56,3,-13,-46,42,-49,28,-8,70,-42,3,2,26,-5,2,-40,-26,44,-6,0,3,-16,-4,10,-9,6,-9,-57,-2,-20,-36,27,-47,-11,-16,-15,-50,8,36,-1,7,-12,-8,3,3,14,-8,15,-7,-1,-27,-2,1,5,1,42,16,18,-6,17,2,-4,-45,3,3,-4,-1,61,-11,-6,41,47,12,9,9,8,-29,-2,27,-6,-17,7,7,0,-21,40,0,4,-4,53,82,-19,3,-20,39,-55,2,-47,-9,-3,-34,-14,-1,-32,-23,0,1,-9,1,22,-37,9,5,-25},
{-37,51,0,-6,-26,-2,-4,-20,0,-28,-9,16,-45,-3,16,25,-8,-49,5,8,-8,-9,6,23,9,36,-9,3,-17,25,-1,16,-2,11,0,-53,-17,4,21,8,-26,5,-4,8,31,0,13,-6,6,17,-5,17,73,12,-5,-3,-5,-8,-4,-52,-3,1,50,29,-10,-33,-7,8,-39,-1,6,8,3,11,36,-36,-34,-24,34,23,4,19,25,-19,-64,4,12,-1,-8,-49,12,-71,13,-4,8,39,-5,31,36,-21,61,-15,-22,-5,4,-4,0,-62,-4,53,-1,1,5,-22,-1,-19,7,55,-20,-13,-4,-11,14,21,23,-1,4,-5,-2,5,11,20,-3,16,-15,-13,-17,5,1,-9,3,-11,37,-7,-1,-13,23,3,-57,-5,26,0,6,68,-6,6,33,47,-7,-8,-12,1,-39,-6,10,5,-20,33,6,-4,-3,49,18,1,5,56,65,0,-3,-5,6,-28,9,-33,-20,-6,-22,1,-6,-21,-13,-32,0,-46,8,39,-47,-22,7,-40},
{-26,38,-3,3,-25,4,5,14,12,-10,5,3,-49,13,3,41,6,0,-11,6,3,-11,-8,14,-8,41,-18,-3,4,28,-6,37,5,14,-8,-35,-7,0,-8,2,-4,9,13,9,-6,-3,-4,0,6,-6,-5,13,67,17,5,-12,6,1,-13,-39,2,-15,1,-15,-10,-31,-21,14,-31,19,1,-15,8,-3,36,-16,-9,-9,-6,50,-4,20,27,-16,-52,-31,3,2,-9,-19,11,-25,-15,3,4,32,13,37,33,-23,22,3,-14,0,-7,3,-21,-1,-27,52,-9,-11,-19,-13,-4,5,6,-2,23,-8,-18,9,-3,40,24,-5,14,-42,11,0,11,35,-1,0,-22,-39,-21,0,-6,1,-6,9,8,-31,0,-22,37,12,-36,-2,5,7,0,18,-11,5,7,42,-9,-5,-3,8,-54,4,-6,8,2,23,13,6,11,36,65,9,0,73,10,-3,0,1,7,-4,-5,0,-13,-10,1,0,-13,-48,-35,-9,-12,5,-8,34,-20,17,-4,-27},
{-29,12,0,34,-35,23,5,37,9,0,0,-31,-2,0,12,-8,11,-3,0,1,1,2,11,7,-17,9,18,0,52,84,5,-28,17,-26,-14,-16,13,5,-49,-31,28,-1,0,17,-50,-38,8,-3,0,-3,-9,-30,33,40,17,-6,37,7,21,-6,30,-20,6,-26,21,10,-2,-3,-22,56,1,-23,-15,-4,30,-5,12,12,-81,37,-2,1,9,-25,-21,-66,0,-7,-31,43,6,-33,-61,-6,13,-5,16,6,18,-26,0,40,-25,14,8,-2,-28,-23,-29,-11,-45,3,54,-8,-3,13,19,-36,56,-6,-33,1,-12,23,10,-5,-29,-3,33,2,0,19,4,-15,9,-7,-7,7,1,3,7,-37,16,-7,-4,-14,34,-3,-26,-10,-47,-3,7,5,-7,-7,16,35,2,-1,11,-2,-40,-2,-1,-6,33,-34,32,-5,14,-10,28,-5,1,86,8,27,6,2,-22,15,-5,42,-19,9,56,30,-13,-26,31,36,-13,49,-9,35,-30,15,10,-61},
{17,-24,-8,-9,-80,-17,-8,50,24,-19,11,-84,22,3,-11,-27,-1,20,-39,-2,6,0,0,18,-25,-2,27,-4,-2,-5,-7,-31,-5,34,15,14,27,-1,7,-46,-31,-6,3,8,-32,-16,27,0,-6,27,0,-43,-14,37,0,-47,39,-4,0,-34,90,8,-13,-21,16,10,3,-9,51,-35,42,-5,18,-4,-20,-6,5,-8,-88,-12,-5,-58,-3,-83,25,2,43,3,-13,36,-25,-16,4,3,33,2,2,-4,34,11,-3,22,-6,19,0,0,-27,-2,-27,-11,-68,-2,0,37,4,-6,14,-28,14,9,-31,20,-24,-16,3,6,11,-15,8,5,11,-34,-2,17,40,17,-3,-10,-2,-5,0,-14,22,-1,-53,-8,-2,-7,-13,-10,6,-4,5,15,20,6,44,-14,-3,17,-1,8,5,-5,1,-4,113,-66,19,69,10,8,-18,1,4,48,-24,7,7,-50,35,20,6,-41,-18,3,-23,-12,15,11,98,24,0,47,0,-17,6,18,-3,-34},
{38,-49,5,-33,-23,9,-6,-13,11,5,-2,-78,-7,-18,-6,-35,3,15,-4,7,3,2,6,29,-27,-7,-14,-3,-59,-81,-3,-7,-15,59,38,41,6,1,54,-17,4,-5,-1,-4,19,42,12,0,8,1,-21,-74,-75,-31,-1,-56,-5,-1,-9,0,31,23,-16,-17,-57,8,0,-19,67,-59,49,-3,0,0,-79,0,25,24,0,-68,-8,-79,31,18,-9,90,38,0,0,62,-25,19,33,0,18,74,-15,-66,16,-13,2,-45,-13,-7,-4,3,51,16,8,2,59,-6,-19,50,0,34,1,7,-27,7,-19,-10,-72,38,-32,0,24,-20,3,-1,10,5,9,66,38,8,-13,3,7,1,6,-13,-16,5,-77,8,10,2,28,-13,11,9,-4,13,7,-8,11,-53,-8,-1,-6,5,5,-8,25,3,34,8,13,-3,-2,-2,-41,6,-5,-34,-25,13,0,0,13,-19,-1,-88,6,15,-70,-14,17,22,-11,-33,6,7,1,-77,20,19,2,-2},
{21,13,-3,-29,34,16,-13,-52,-11,-3,-4,30,16,17,0,-25,-4,-27,-13,2,2,12,1,25,-15,-1,-54,-4,-71,-58,0,3,29,12,4,35,-37,1,-9,31,36,-4,4,-22,25,-1,1,-3,2,-36,-1,-119,-44,-25,-14,1,-50,2,-25,-6,-39,-91,-15,5,-67,8,0,24,18,-23,5,-7,-34,2,8,-9,-1,14,12,-58,3,-100,29,32,-1,92,32,-12,-8,81,-9,14,45,5,-15,57,-1,-1,-26,-18,19,-64,3,5,0,3,53,11,25,-5,105,-1,-13,55,-3,39,58,22,-37,-3,7,-1,5,14,-43,-6,26,14,-20,-6,-8,4,-4,41,-5,15,12,-12,-4,-3,-2,10,-20,-1,-15,11,2,6,20,3,-9,-67,0,16,-35,7,2,-30,9,-6,-1,0,-42,5,-13,0,-49,30,-6,-64,4,-3,-31,-5,4,0,-4,1,2,34,-8,-25,-3,-50,14,0,-86,15,-7,0,-140,-22,-3,3,2,-81,21,17,-3,11},
{-3,14,-1,-21,22,17,-10,-19,-69,-49,-1,56,7,12,11,-16,4,-51,-12,6,0,1,10,29,27,-1,-45,-1,-38,-7,0,22,40,-21,-19,9,-46,7,-21,26,40,0,14,-35,7,-40,0,-2,6,-41,5,-107,-24,-32,-42,33,-53,-7,-56,-10,-60,-107,-2,21,-98,5,-2,38,-40,-5,-19,3,-27,-10,-2,-13,-30,-3,4,-37,-2,-95,29,21,-7,33,12,5,-4,10,25,-15,30,-2,-34,6,-3,25,-76,-27,18,-33,-30,31,-2,-4,29,20,0,-21,70,8,9,38,-12,21,12,68,-29,-4,-3,-21,26,-3,-36,2,-3,3,-29,-2,0,2,0,13,-33,18,26,-8,-2,3,4,13,-13,0,11,-8,57,-6,11,7,-11,-94,5,1,-15,-8,-4,19,12,-16,-12,8,-89,3,-36,5,-70,33,-12,-21,-4,-10,-1,-8,0,50,20,-35,-9,45,21,0,5,-22,6,1,-83,67,-81,-3,-81,8,-1,23,3,-27,36,24,5,22},
{-42,-6,-8,-3,2,-6,2,22,-44,-75,-4,15,14,-10,-28,29,-5,-14,15,6,-2,2,-5,-10,30,-15,-60,-11,-51,38,-3,1,-17,10,-27,15,-21,-15,-3,4,17,-4,-9,-50,3,-25,-5,0,-1,-29,-7,4,-20,-16,-36,16,-8,-3,-15,-2,-50,2,0,-22,-72,-18,-29,-36,-30,-15,-11,-28,-8,-3,-11,2,-10,-22,-5,-47,-3,-69,-5,-4,-109,23,11,6,17,-65,16,35,9,0,-77,38,-15,22,-13,-80,-31,-21,-25,-47,-3,-1,-7,-4,-31,15,-8,-16,-25,0,5,1,-71,-32,38,-18,-5,-5,27,17,3,0,-21,-23,-13,5,-5,6,-4,33,-36,0,18,-3,-8,3,-8,-6,-9,0,19,12,19,-22,-56,-31,16,11,4,-3,-7,-8,1,25,-20,-22,-2,2,-24,5,-34,7,40,26,16,-55,21,3,30,1,4,14,14,-6,-9,-5,-23,6,4,-23,1,-2,-122,34,-119,10,-24,11,-18,3,7,7,2,-43,-4,-33},
{-11,29,8,-22,-123,-15,-7,-11,-7,15,-2,-3,23,15,-42,-26,-12,-19,-18,-2,0,-3,-9,-21,-19,-54,-3,0,14,-29,-5,-59,-25,-6,-11,11,14,-36,-96,-13,-21,0,24,0,-16,-19,-70,0,5,-22,-32,-19,-41,-43,-6,-11,-35,0,-32,-1,-11,29,-52,-4,-18,0,-10,10,-5,-12,-36,-22,-45,3,1,-26,22,-18,0,-26,2,2,-3,-43,-19,-13,-13,3,-9,1,-38,30,1,4,-40,-26,-28,4,24,9,14,-4,-23,-28,-5,-4,-3,7,-21,-17,-11,3,-34,-27,0,1,-61,24,-12,-30,-18,-7,4,-23,-15,-1,-56,7,-17,-9,-1,-239,1,-13,3,2,20,-8,3,-2,-7,7,-11,3,-10,-13,-26,-25,15,10,-23,5,7,-53,-20,-1,5,-29,-32,-8,13,0,-10,3,-6,8,6,-6,-8,7,13,-14,-8,0,1,-44,-21,8,-10,-14,-4,25,1,-23,-5,-8,-11,18,7,44,-6,0,-20,3,2,-6,14,-24,-8,24},
{43,37,-8,-35,-10,-12,-15,24,-15,21,-10,2,14,34,16,-151,-9,-22,24,8,4,-8,-10,11,-21,-30,12,0,41,-116,-9,-14,-20,-8,-5,17,16,11,12,-1,-55,-2,25,-14,-7,-82,-56,-3,-4,-11,-57,-50,-41,-26,-17,-2,-35,-1,-5,-44,-33,-65,-20,23,-19,-7,-8,19,-23,-60,-55,-13,-44,-9,63,-31,45,24,-10,-67,6,-44,3,16,-52,-55,14,-8,-64,52,-64,188,19,1,-1,36,-14,-24,33,-7,22,44,7,-96,-6,-10,12,10,-23,-20,-14,-4,-16,0,6,49,-115,56,-4,-23,-21,-13,41,21,-12,1,4,3,-22,-1,-1,-41,-6,-56,-7,-6,17,-10,2,1,-1,43,-27,0,0,-22,-23,-1,22,1,-47,0,1,-24,-7,-1,11,18,-45,-41,34,2,-37,-7,13,3,-30,-11,-8,3,-1,-33,-3,0,-3,-13,-84,21,-7,-37,-21,39,-12,9,-12,-50,16,-20,19,6,22,28,-3,22,-3,-22,6,-44,1,38},
{17,27,4,-25,-15,23,2,16,4,4,8,12,28,12,34,-87,-2,-4,-11,-2,-6,12,-3,46,-11,-22,12,-4,21,-39,-8,3,-16,-17,-1,2,25,5,17,5,-8,-4,-18,0,-15,-93,-17,6,0,4,-57,-96,-3,-22,-39,39,11,-10,-20,-49,-104,-128,-62,31,-10,-39,-3,11,-25,-55,-65,-4,-10,-1,9,-14,-79,-63,-74,-66,-2,-105,18,0,-58,-31,45,7,-70,76,-17,70,83,0,-21,71,0,12,5,-24,48,28,-24,-110,-2,0,0,24,39,18,15,-9,-28,57,-4,104,-57,40,-33,-6,-16,-8,27,24,-47,-1,41,-33,-10,-2,-7,-21,-2,6,-23,22,53,-7,4,6,-3,24,-46,-34,25,-38,-15,9,36,-10,-31,-18,2,-16,-17,-1,25,8,-29,-23,5,2,-78,-8,16,0,-58,-44,21,-18,-31,-42,-20,-7,0,-15,-106,11,-4,-49,6,60,-9,17,-4,-46,33,3,31,12,11,7,-4,42,-7,-39,31,-3,4,57},
{-11,13,7,-18,1,-7,-3,9,26,20,10,5,2,9,39,-48,-2,-2,-96,5,3,-8,3,52,-35,-7,-37,0,2,25,2,-31,-9,14,-1,-2,37,14,-2,-17,53,-3,-25,0,2,-48,31,-5,1,-23,-3,-120,34,-10,-19,49,21,4,-22,-28,-77,-69,-27,39,-18,-3,-12,20,-13,1,-26,0,-28,-2,-46,12,-85,-25,-24,-28,-7,-134,-32,22,-76,-17,28,0,-10,67,-29,12,30,5,-51,85,-14,-4,-5,4,26,-20,-6,-61,-6,4,7,10,31,17,23,8,-2,63,3,81,-50,-13,34,-8,20,7,-3,15,-106,-4,31,-16,-17,3,5,19,-7,-3,-5,-8,64,3,3,2,3,9,-45,-44,14,8,-14,-6,32,11,-26,-4,1,-8,-69,3,30,-9,-24,-34,-23,-3,-65,-1,31,7,-37,-7,22,-101,-11,-35,-59,5,6,-24,-46,1,3,-5,9,43,2,-18,17,-46,-32,6,9,16,15,-4,6,49,0,-34,43,26,-3,5},
{-85,-21,-7,-18,54,-40,13,3,26,2,-1,-6,-41,-2,47,-37,3,44,-40,5,1,0,4,40,-31,24,0,-7,-38,72,0,-35,-19,22,8,-22,35,5,-7,6,30,5,-35,1,-12,3,-25,0,8,-6,22,-31,58,7,24,-3,-13,6,0,27,30,4,15,34,-43,2,-26,-48,6,-16,-32,-8,1,-13,-39,38,-50,14,1,-25,-4,-112,-33,6,-4,19,37,0,30,40,-29,-48,27,6,-30,16,-3,-11,11,14,-15,-69,1,-30,-2,9,35,14,18,44,22,0,16,22,-4,44,-43,34,22,-8,13,15,-9,-5,1,0,29,10,-48,7,-2,17,10,-39,-20,-11,65,-5,5,-2,-5,29,-18,-1,-30,32,13,0,-23,31,-27,-27,2,-5,-19,-2,16,-11,23,-24,-82,6,-15,-2,29,3,-54,88,23,-59,-18,-9,-30,4,0,-5,38,-66,0,13,22,-4,-7,-25,16,5,-77,-12,-12,-9,10,-3,-8,29,6,0,-16,1,2,20},
{-76,-22,2,-37,25,8,10,-37,5,6,-5,15,-21,-21,20,-13,5,-17,16,0,-5,-8,0,32,-7,52,11,-9,-37,65,0,-3,-14,21,-11,0,16,-1,4,33,-6,-9,-25,-6,0,-6,1,2,-6,-5,-23,29,65,23,38,-30,-8,-3,27,17,94,70,49,24,-34,-16,-26,-1,-33,-8,-23,-29,-18,2,13,-21,-25,-2,31,0,-3,2,38,-7,-8,13,20,5,6,-38,2,-81,33,-3,37,-1,-4,5,15,-24,7,-78,-34,37,-7,-2,7,-8,-11,35,40,11,2,-14,1,10,-3,39,8,-21,-30,-2,-21,-7,39,8,17,-1,-20,-3,2,21,0,-5,-28,-32,-1,0,1,5,3,7,32,25,-39,-10,0,0,-61,-24,10,-38,5,21,-3,1,54,18,40,9,-46,2,-13,0,35,0,-13,34,8,4,0,27,11,4,0,7,66,-41,-6,1,36,-22,0,-16,2,-6,0,25,-35,-21,-5,12,0,15,10,41,-39,-37,1,-1},
{-31,9,7,5,-2,4,-9,-16,9,-9,11,49,-41,-6,-9,14,2,-60,0,6,1,-2,-11,6,-11,55,-19,0,-2,43,6,15,-20,1,-9,-20,-45,-8,-1,1,0,-7,39,7,9,-5,20,9,-7,-9,-3,29,75,-17,14,-19,-6,-2,-15,-58,-3,67,16,-3,-6,-25,-25,24,-37,5,0,-49,-5,-4,-3,-36,-20,-55,23,22,-1,14,9,-10,-20,-9,-32,-1,2,-21,1,5,20,-9,-35,41,10,16,42,-14,44,-25,-54,-19,1,-4,-38,-67,-38,20,4,4,-50,-9,8,7,-11,48,4,-45,-4,11,-34,40,14,-2,25,-1,-5,-9,5,26,4,15,8,-27,22,-12,0,-6,7,8,40,-24,1,-19,9,-1,-45,-8,34,13,2,11,8,-10,83,37,-11,11,-2,-8,-33,2,6,1,-12,-4,0,6,6,49,81,4,1,31,30,11,1,6,38,-9,-3,-16,13,-4,-15,27,-9,-17,-7,-19,5,-5,6,46,-3,-41,8,-43},
{-13,-2,-4,-8,-25,-4,-12,49,-2,-19,2,15,-49,22,8,1,3,22,7,-7,-7,3,-10,-4,-2,21,-12,-8,36,33,-3,-16,15,11,-26,20,-1,26,-19,-19,34,4,49,14,-27,21,-15,-4,4,0,-2,-20,55,21,23,-30,-13,6,2,-29,-9,-41,-2,-38,-8,-33,-20,-8,-32,8,-8,0,-6,-2,36,-13,5,-2,-25,35,-5,-1,13,-19,-13,-63,-6,1,35,-20,-18,-89,13,4,8,20,5,8,39,-25,-24,18,-16,-30,1,0,-56,0,-34,2,-48,6,-49,2,7,43,18,-27,25,-6,-15,13,-28,48,7,-7,-41,-20,8,5,0,48,-3,9,-18,-13,-18,-1,2,8,4,64,30,-6,7,-34,6,5,-35,-9,6,0,10,-26,3,-6,25,42,-18,-11,7,-3,-11,-8,-41,-3,-3,30,-15,15,13,10,48,5,7,63,-12,8,-5,12,2,22,-5,57,1,-10,-31,52,-12,-34,9,21,1,22,6,14,26,3,-5,-48},
{-14,-8,2,22,-55,14,11,68,-13,4,3,-87,-14,16,29,-27,0,20,-2,5,-5,-4,-2,0,-43,-11,24,1,38,36,-4,-47,51,-21,-34,42,33,11,-57,-24,24,5,-2,4,-69,3,-9,-3,6,-33,-11,-45,70,57,48,-20,4,-2,45,-7,55,39,-5,-26,57,8,-29,-27,-39,37,7,-32,7,3,32,-15,5,15,-46,29,0,3,-28,-6,26,-73,5,-4,37,1,-44,-124,-84,0,18,17,9,-9,19,-18,-36,46,1,-4,-7,4,-37,7,-35,13,-77,0,18,2,1,22,50,-30,56,8,-17,10,4,1,-6,8,-14,18,2,2,5,3,6,14,-1,4,-8,0,-4,6,-2,-3,8,2,13,-35,13,-8,-52,-3,-26,-10,-2,-6,11,8,2,23,-7,-22,22,0,-10,-8,-20,-5,26,18,38,9,22,-8,28,9,-8,47,-18,13,0,36,9,22,-3,80,-46,19,-47,63,-3,-24,61,84,2,60,-7,28,-37,10,10,-85},
{-9,-50,1,-26,-40,-8,-22,63,-2,-28,0,-153,-7,-8,0,-5,0,28,-48,-3,9,-3,11,20,-19,-7,35,4,19,-49,-3,-7,-3,7,-25,9,40,13,34,-13,-30,8,11,-7,-31,27,37,-5,1,44,6,-4,70,37,6,-41,36,-5,-3,-33,72,115,-5,-16,13,-1,-21,-21,-11,-28,47,0,5,-2,-49,-20,11,-52,-70,1,-7,-55,-7,1,11,-12,-13,-6,3,0,-37,-56,-56,-7,33,20,4,-11,19,-9,-28,7,0,9,-3,1,-8,54,-15,-1,-52,2,3,29,3,-43,7,11,62,2,-34,13,-12,-40,14,-4,27,-16,24,7,4,-64,0,110,37,-15,8,0,9,2,-1,-17,15,-19,-31,-37,6,2,-22,1,66,37,8,0,20,6,18,-3,0,1,-35,0,12,8,-22,3,102,-29,-40,98,36,13,3,5,5,-20,-53,8,0,14,39,-10,0,-9,-13,-10,-70,-25,41,6,101,43,0,41,2,29,-12,13,1,-36},
{13,-50,-7,-69,4,0,12,-29,1,16,1,-44,0,-39,-5,-33,1,26,-31,-2,-6,5,8,26,7,-4,-28,0,-10,-100,0,23,7,24,11,25,-21,17,19,25,-18,0,-2,-1,46,42,13,-2,2,28,-20,-2,-20,-5,-9,-17,8,8,-19,-5,41,-43,-49,-14,-40,9,-14,11,1,-86,33,18,-5,9,-92,-31,38,18,-7,-59,-8,-52,14,19,-14,29,10,-6,-32,25,-13,-27,-3,1,40,33,-11,-55,-5,27,16,-74,23,-21,5,8,11,38,10,29,64,-9,-14,30,7,-19,14,11,8,18,7,-26,-59,10,-47,1,24,-7,13,9,-1,-5,-4,102,24,-21,22,10,-3,-2,0,-41,-12,-10,-20,-29,17,3,17,21,29,8,0,29,-33,3,-7,6,16,26,-23,-4,-6,5,3,1,3,-9,-6,38,30,5,-19,3,8,-39,-53,11,7,22,2,-18,-4,-67,15,-13,-72,5,50,9,8,-46,1,13,0,-39,-3,3,0,30},
{24,0,-5,-51,35,10,-1,-66,-23,19,-3,39,2,18,18,-48,-5,-28,-17,-4,1,0,-3,29,24,5,-47,9,-24,-37,2,19,62,-3,9,21,-58,14,-40,29,24,0,11,-22,38,-24,0,-7,-9,-13,2,-32,-38,-23,-11,25,-52,-1,-28,0,-35,-139,-29,-16,-58,17,-12,48,-25,-47,-5,20,-35,3,-26,-28,21,0,12,-106,2,-81,23,12,-26,27,-1,6,-10,30,19,-23,41,3,23,24,-5,-22,-37,24,18,-88,19,-20,7,3,13,22,13,7,87,12,14,25,5,6,105,20,-19,10,28,-17,-16,1,-36,-2,12,13,-7,-5,1,0,0,41,-1,-14,13,-10,5,0,6,13,-10,1,-3,-8,11,1,26,22,10,-67,6,17,-30,-2,-11,26,25,10,3,-4,-38,-4,7,5,-63,8,-25,-31,11,-4,-33,5,7,-17,-2,-3,0,28,10,-16,8,-54,30,-4,-74,57,11,4,-155,-23,-6,4,-5,-36,-1,6,-2,18},
{39,2,-4,-35,10,12,-15,-32,-48,-46,0,49,6,2,-11,-1,16,-31,-16,0,-7,-2,-6,25,49,1,-61,4,-11,-13,0,12,57,-23,-12,15,-65,12,-35,23,12,-4,7,-51,3,-47,-10,-4,-1,-13,13,-38,-13,2,-66,38,-36,4,-22,-18,-37,-142,-11,19,-125,6,-20,32,-59,-28,-19,0,-26,-1,-13,-18,-14,0,8,-85,-2,-70,10,-8,-34,-12,-10,-6,22,-62,22,-10,17,3,1,-24,-22,4,-81,-2,27,-67,-10,-16,5,4,13,20,-6,0,53,7,15,10,-9,15,35,46,-21,10,13,-15,27,-18,13,-4,0,9,-10,-10,4,5,0,1,-11,5,15,7,0,0,-1,8,-10,2,1,0,25,-20,8,18,-12,-99,3,14,-15,-2,-13,58,2,-3,-6,-2,-64,-2,-1,0,-45,13,-19,2,10,-1,-26,4,6,26,26,-22,-9,25,14,0,-2,-11,12,5,-63,65,-56,13,-99,-17,5,21,-4,-8,6,6,0,24},
{-12,-21,6,-20,0,-12,-5,-21,-34,-42,-6,10,-75,-11,-44,16,-15,-5,-3,8,3,-9,-8,-5,24,7,5,-1,-17,12,6,-6,23,-4,-20,18,-42,-7,-13,-1,-1,-5,-1,-32,-9,-7,-5,1,-6,-7,-15,11,14,11,-5,10,-14,-1,-2,-33,-30,66,-30,-27,-60,-18,-27,1,-49,-51,-21,-10,-13,1,-82,-10,9,-35,0,-50,0,-20,-6,1,-147,8,-14,7,23,-84,4,15,-2,-2,-42,10,-11,52,-29,-26,-19,-36,-9,-26,3,-6,-5,-6,-54,0,-21,11,-11,-14,-11,0,9,13,44,-22,0,-9,34,20,0,-5,-10,-6,-7,-2,-1,19,0,13,-11,7,5,2,-3,-4,-1,-21,-9,1,4,-1,3,-8,-164,-17,4,-14,6,0,-5,3,-9,17,5,-15,-14,-7,-23,-1,-22,-6,29,23,-11,-19,17,-8,33,-5,-8,11,5,-4,2,12,17,-4,-2,29,1,-9,-76,-44,-85,-25,-8,12,-14,-18,-9,-9,-15,-12,0,-12},
{-44,29,-7,-1,-44,-16,-17,16,16,3,4,7,14,22,-31,-75,-12,-7,2,-4,-2,-3,3,-31,-23,-44,-9,8,25,-94,-5,-25,-38,-18,-5,-4,14,-29,-55,-3,-24,0,21,0,-8,-26,-44,-1,-2,-9,-20,-20,-40,-26,-8,-13,-27,-4,-22,14,-53,50,-36,6,-31,-21,18,8,-10,-4,-63,-8,-55,6,54,-24,40,-26,-3,-27,7,-25,-2,-73,-205,-24,-20,-5,-12,10,-42,-62,18,6,-44,-55,-13,7,24,2,9,33,-2,-104,-6,6,-8,-15,-132,-20,0,-10,-39,-23,-5,14,-113,2,11,-34,0,3,-7,-10,-7,2,-24,18,-20,-4,-1,-36,6,-7,-6,9,-1,0,-2,-4,4,25,-21,11,4,-9,-38,-11,-6,12,-21,18,-8,-34,-22,-1,-11,-30,-55,-26,11,-2,-10,0,-16,-8,11,1,-19,-4,2,-26,-31,7,7,-21,-57,18,2,-9,0,0,6,-11,-23,-15,-12,0,3,5,5,13,-22,-4,0,8,33,-37,0,30},
{72,52,7,-20,-19,-6,-21,23,-7,5,-3,-7,9,32,15,-117,-8,-6,25,1,-8,-5,-9,8,-19,-55,-4,-2,40,-107,-6,-14,-19,-17,0,11,37,7,22,-1,-28,0,23,-6,-2,-60,-25,-2,-9,-10,-36,-40,-42,-33,-20,8,-22,5,-2,-45,-33,-27,-34,21,-20,-5,6,6,-30,-62,-107,1,-31,-2,71,-8,15,48,-15,-133,-3,-44,0,9,-59,-57,-2,2,-55,48,-40,137,50,-10,-14,34,-13,-5,30,-22,23,98,5,-258,1,-6,6,10,-30,-15,-7,-7,-41,-25,8,-60,-90,33,-1,-18,0,-11,9,24,22,5,-14,5,-6,1,-6,-32,6,-60,0,-7,11,-6,6,1,-3,48,-18,-4,-2,-21,-8,-4,17,-3,-32,14,7,-19,-4,-3,-3,21,-71,-29,17,-4,-35,0,13,-2,-43,0,-20,-10,1,-31,-12,-8,7,-16,-92,22,3,-36,-21,24,-12,4,-2,-43,1,-13,10,17,22,19,7,6,-5,-18,10,-47,-1,49},
{59,16,0,-10,-55,32,-14,12,10,-7,-1,28,26,46,15,-76,-9,-8,17,-2,-1,12,-4,18,8,-32,11,-1,46,-64,-3,-22,-20,-13,10,9,17,23,29,6,-7,-3,29,-8,-10,-79,-30,-4,0,16,-70,-52,-13,-7,-20,24,10,-5,-7,-47,-61,-122,-65,34,-11,-26,-3,9,-21,-47,-73,2,-3,2,5,-6,-157,34,-18,-87,-7,-79,35,8,-35,-50,12,-9,-53,52,-25,114,56,5,5,51,5,-7,7,-29,43,18,-22,-315,0,3,-7,23,18,-2,20,-14,-36,11,-3,74,-43,24,1,-2,-21,-9,6,28,-37,4,12,-37,0,1,-6,-5,-1,2,-10,10,34,3,7,-6,-7,49,-38,-33,19,-62,-1,2,20,-12,-5,-7,-1,2,-13,-3,-11,21,-97,-7,9,-8,-49,7,16,-2,-63,6,8,-2,2,-53,-21,7,6,-40,-105,31,1,-50,1,52,-2,18,5,-53,3,-13,3,14,15,8,9,1,0,-34,20,-2,0,39},
{37,10,-1,-19,-36,12,-17,0,10,5,1,3,20,27,17,-41,-2,9,-61,-2,-4,4,6,29,7,-18,-25,-6,52,-8,-4,24,-8,7,0,11,26,21,42,-41,14,5,-3,-2,-32,-65,10,-4,9,16,-20,-91,11,11,-19,51,14,-6,-2,-40,-32,-83,-21,59,-13,-18,-7,14,-15,-30,-49,7,-4,3,-28,9,-84,44,-16,-66,-8,-101,0,-1,-57,-41,20,-10,-20,14,-26,57,45,-8,17,88,-26,-14,18,4,32,-28,-1,-170,2,-8,4,1,16,-1,44,-2,5,28,2,82,-4,-67,-7,0,-1,-17,-7,33,-79,3,28,-20,-18,-4,-4,14,-2,-25,-6,9,42,-10,2,-5,0,40,-80,-51,-6,-23,-2,-6,35,4,-5,-27,6,-8,-35,0,0,-16,-66,-4,1,0,-35,-5,42,1,-36,-6,26,-68,2,-68,-34,2,1,-85,-107,32,1,-54,-27,68,4,20,26,-52,-43,-1,-14,36,19,-9,-4,11,-3,-23,20,23,-2,-2},
{-17,-38,-2,-74,32,-46,-11,-9,-20,7,8,-10,7,1,37,-32,1,35,-55,-2,9,10,12,50,-11,28,-6,-1,45,60,-2,27,8,25,-4,30,31,22,-6,-17,26,5,-33,-12,-19,-29,-13,-7,-5,0,-8,-57,34,50,19,27,10,4,22,-39,5,-21,34,39,-21,4,-37,-35,13,-37,-66,-8,-32,7,-51,7,-28,36,-10,-9,-5,-99,-27,6,-28,-25,4,0,17,-1,-32,48,32,-1,-33,47,-11,-13,21,7,-1,-55,7,-64,-4,7,10,0,-6,23,54,11,23,14,2,52,1,-37,22,-4,1,4,-8,-39,-44,9,19,21,-13,-7,10,18,5,-78,10,-12,56,3,3,-8,-4,3,-85,-4,-12,21,-9,-12,14,12,-43,-35,2,-6,-35,9,1,-36,6,-18,-58,-8,1,5,57,4,-54,43,32,-39,3,-79,-22,0,-2,-74,-51,-21,-5,-30,-44,41,4,17,34,-13,-37,9,-37,38,11,4,10,4,-2,-40,-16,-63,-6,27},
{-43,16,0,-63,-11,-9,-11,-38,-19,6,6,7,16,-14,19,3,11,5,14,1,-3,13,5,48,-24,32,1,-7,12,57,3,10,-9,9,2,21,11,6,-19,6,31,-5,-13,-4,-12,8,-15,9,2,-17,-30,-16,45,27,60,-12,-9,0,-9,-89,56,102,28,9,-26,-6,-48,-9,21,-34,8,-38,-6,0,-14,-48,11,-22,25,16,-5,-47,12,30,7,21,-6,0,30,-7,-41,33,10,-9,-53,39,-3,10,8,-19,23,-43,-58,34,2,1,-34,-82,-62,14,28,-4,4,-5,0,54,-26,58,-1,-39,-36,4,11,-3,0,-1,8,4,-38,1,-4,27,4,-34,15,-11,37,-10,10,9,-5,-10,-24,3,-24,-35,-18,-11,-1,-46,0,-24,9,14,-3,12,-8,17,57,3,-58,-5,22,0,28,0,-75,67,22,8,26,-28,59,8,-4,-65,-40,-33,2,-26,16,49,0,-5,22,16,20,61,-37,9,-38,-3,5,7,7,21,-21,-76,-6,22},
{-15,20,8,-10,35,10,-1,28,4,-29,7,26,5,24,-7,12,1,-16,-13,6,1,2,-4,2,-7,29,-41,3,18,9,10,-56,24,-2,-11,-5,-38,19,-5,5,5,5,67,-12,-21,36,-15,7,6,13,5,-6,39,27,20,-39,-30,0,-28,-88,-11,-13,-28,-14,-24,-7,-40,-19,26,-20,-8,-31,-7,0,-61,-12,6,-33,-27,4,7,6,-5,41,46,5,9,0,46,-31,-31,0,31,-3,55,31,0,-17,9,-9,8,4,-55,-16,-5,-1,-41,-38,-64,-3,-46,8,-73,-17,-2,51,-4,67,29,-28,-19,-17,-7,32,42,0,-43,-31,-9,-2,-3,26,-5,0,41,-15,40,0,2,1,1,96,57,0,-7,-27,-10,14,-5,-38,32,22,1,-2,20,0,66,42,-19,13,-30,4,69,-7,-42,3,-16,6,-33,-14,41,-29,60,3,1,-60,-12,-3,7,-8,23,45,-4,1,28,20,-18,39,2,-29,-2,2,11,24,-6,16,11,-30,4,-32},
{-27,13,3,-14,3,10,-7,62,-1,10,10,-1,5,33,-4,-30,0,15,13,-4,-6,-2,5,-19,14,-31,-54,4,0,-44,9,-32,67,2,-8,59,6,1,-14,-33,7,-5,15,-7,-32,52,-22,6,-1,11,-13,-10,21,41,25,-42,-30,1,29,-25,11,-46,8,-18,-27,-10,-34,-35,11,-2,9,-12,5,-2,-53,17,9,34,-53,12,-8,25,6,62,84,15,37,-1,49,-41,-61,-156,28,12,119,23,6,-43,10,-26,-77,44,-3,-38,5,-3,-27,39,-67,-39,-43,0,-14,11,3,59,66,-6,11,-5,-13,-3,22,-8,22,9,0,-7,-21,5,0,33,-5,5,-49,22,-37,-3,-4,7,-2,115,38,8,-29,-33,-2,1,-6,-20,-28,-6,-5,-17,7,-9,22,38,-5,-19,1,-1,56,4,-41,-1,12,53,-42,1,25,-20,1,-5,-7,3,17,14,0,17,28,40,-5,68,-38,-3,-50,6,14,-33,49,50,11,-6,-7,-8,21,24,0,-49},
{-15,-47,-7,14,-13,20,-1,49,-11,-3,2,-104,9,12,18,-9,0,1,-8,8,-7,11,2,-8,-26,-62,24,1,8,-23,0,-58,50,-29,-34,54,45,6,-9,-7,-31,-8,-3,-14,-32,43,44,0,-6,-18,-5,-7,60,24,28,-22,-8,5,29,-5,5,96,32,-9,1,-1,-16,-11,-24,19,15,-55,23,9,-22,-8,-10,-29,-10,6,3,38,-14,63,68,17,16,0,21,-31,-51,-120,-95,-9,-2,-11,3,-36,-43,-9,-75,20,11,-3,-8,0,22,41,-4,-22,-11,4,27,-3,-10,25,47,4,33,-12,7,0,50,-58,-7,7,54,4,10,-8,5,-34,7,20,-15,39,-32,9,-1,9,7,-30,5,-14,-1,-46,4,10,-2,21,0,14,2,-8,24,-1,10,-1,-2,-32,8,-6,36,2,-24,-8,-10,2,17,40,17,21,30,1,-5,-16,1,30,-4,45,35,5,1,79,-51,-19,-11,15,46,-5,38,90,5,37,-2,33,-43,-1,2,-73},
{10,-55,4,-27,0,-12,9,-9,8,3,-2,-121,10,-6,-17,4,1,0,-33,-6,1,11,7,34,-13,-10,-2,0,0,-78,2,24,0,-21,-7,-9,5,8,58,20,-60,6,-9,0,25,11,33,-2,1,11,-3,59,52,6,10,-15,19,-5,9,-16,26,42,-15,10,-8,15,1,16,-39,-23,28,7,-2,5,-55,-21,1,-51,11,32,0,0,-8,50,28,30,-15,-8,-14,-45,-56,-165,-87,-3,-2,-14,11,-8,-43,18,-1,-35,11,26,6,3,-5,38,-2,11,58,10,3,15,4,-65,21,30,75,14,-8,17,36,-42,1,7,55,1,1,0,-12,-69,5,41,11,-20,7,2,0,-8,-2,-43,10,-39,18,-44,-24,12,12,29,57,39,-2,9,0,-8,15,14,25,0,-24,5,43,2,-7,-3,-2,-32,-26,78,16,10,17,-4,5,-56,-49,11,0,6,28,-6,4,9,-9,-37,-7,-44,60,8,20,-30,-5,-8,1,34,-53,24,4,-9},
{27,0,7,-72,21,-8,-9,-67,13,17,-1,20,9,-8,-28,-5,-4,13,-27,0,5,-3,6,24,9,6,-37,-3,-12,-84,-1,23,50,2,31,-13,-55,6,-27,26,-40,0,6,-6,57,35,-1,6,4,-1,-3,68,-6,-22,-30,-14,-7,-6,-2,2,7,-100,-42,-5,-63,21,12,55,-40,-92,0,38,-26,-4,-51,-44,24,14,19,-4,-1,20,17,21,-20,38,0,0,-44,-23,-12,-60,-47,-9,23,-18,4,-49,-36,37,26,-72,28,-3,-5,-4,-18,20,7,29,72,6,9,13,-1,-72,27,35,9,29,19,-22,-27,-6,-21,-6,6,12,16,9,-11,-19,-2,26,17,-40,25,12,-1,2,-2,-35,1,-11,-11,-26,1,-7,26,25,44,-31,3,24,-45,0,2,37,23,16,-21,4,17,2,20,-3,-85,-25,-21,7,10,15,20,-9,5,-48,-46,0,-1,1,16,4,1,9,21,-24,10,-14,53,1,-64,-80,0,-4,0,30,-40,-3,-3,22},
{32,-1,4,-45,24,-10,-24,-85,-10,28,-7,49,-4,4,-3,7,2,-40,-3,-8,-1,-7,0,20,21,18,-25,0,4,-73,2,25,94,-9,32,-2,-77,11,-52,13,-10,5,20,-15,45,0,-17,-5,7,0,11,43,-33,-11,-36,-1,-49,-8,-9,1,-51,-112,-37,11,-88,17,8,50,-59,-26,-30,37,-40,1,-27,-18,6,3,26,-68,0,-9,15,-9,-47,30,-17,-5,-27,-42,19,-28,4,-7,34,15,0,-22,-68,47,44,-70,21,-3,0,-2,-17,4,-2,39,49,-3,13,10,0,-48,99,56,-8,28,24,-27,-23,-23,31,-5,8,25,26,6,4,2,4,-13,14,-31,11,6,5,3,-7,-7,-4,-4,-17,-1,-1,-18,16,18,17,-106,1,22,-32,-2,-14,66,6,10,-5,0,-17,6,37,-8,-122,-12,-25,-16,8,10,-12,0,5,-9,-12,-28,6,19,17,16,6,21,24,-10,-11,0,6,-9,-190,-49,-12,3,3,-6,-30,6,0,37},
{35,-12,1,-36,12,-9,-16,-63,10,-25,7,12,-6,-12,-15,23,-14,-43,-15,9,3,-9,1,9,25,20,17,5,-6,-2,-6,4,69,6,22,-2,-30,-2,-22,0,2,-6,-6,-18,5,-7,-23,-9,-8,-2,0,13,-22,2,-5,19,-44,-9,-14,-12,-20,-65,-17,1,-122,10,0,8,-51,-9,-23,17,-23,-1,-54,-1,-17,-18,16,-113,3,-32,-2,-35,-79,22,-12,1,0,-110,2,-10,15,-5,19,3,-9,-30,-93,27,47,-58,-10,-13,-8,-8,-11,-8,-29,-4,5,-6,14,1,3,2,18,63,-9,6,6,-21,-6,-38,19,-4,-10,0,17,-3,-7,14,6,-27,13,-18,17,-8,-9,0,-7,16,-12,12,-56,11,5,-8,3,4,-13,-54,-9,14,-12,-15,-9,44,2,-8,-13,-1,-28,6,34,3,-111,5,-7,-16,4,2,-1,-8,3,-17,31,-10,-2,25,37,20,-3,21,18,-3,-13,23,-37,15,-72,-38,-19,8,-4,5,-17,11,6,39},
{-29,-43,4,-6,1,-10,-8,-29,-18,-33,0,6,10,-30,-26,29,-15,-14,-1,8,1,0,2,-12,29,-1,-57,6,-34,28,-8,-18,24,8,-15,0,-17,-21,-9,1,0,3,-12,-78,-8,-11,-2,-4,-3,-10,-3,18,11,6,24,40,-12,6,1,-1,16,88,-17,-7,-54,-20,-15,-26,-20,-60,-16,-8,9,-3,-58,8,25,-29,-5,-50,2,-16,0,-11,-88,-2,1,6,6,-59,8,-679,-30,-7,3,-307,-18,17,-23,-19,-17,-60,-26,-30,0,6,-39,-12,-103,-21,-36,11,-7,-17,-6,-26,10,-3,52,-39,-4,11,45,3,-6,0,-17,0,-13,-2,0,23,0,6,0,-2,16,0,1,5,2,-47,1,1,-16,2,2,-16,-43,1,25,-10,0,-16,-10,-10,-20,14,-4,-17,-21,-6,-12,8,-5,5,14,25,5,-1,8,-8,25,-1,8,4,-6,-27,-7,-6,26,-3,7,50,-9,2,-31,-15,-104,31,9,1,-24,-27,-7,-18,-22,2,2,-19},
{-31,11,0,-11,-216,-2,5,-19,-7,-18,-3,4,-29,6,-49,-20,-2,-26,-13,-2,-1,-1,6,-14,1,-1283,-40,5,7,-5,7,-28,-12,-13,2,-2,5,-71,-37,-1,-1,-6,2,-97,-5,1,-23,-2,-3,-7,9,8,-10,-184,-21,4,-28,1,-100,-205,-8,1,-353,-9,-48,-26,1,-9,-6,-51,-85,-12,-16,4,-2,-23,0,-7,-10,-10,0,6,-5,-55,-41,-4,-15,-1,-16,-5,-17,-244,-9,-1,-207,-164,-7,5,26,4,9,-1,-47,-354,6,1,0,-1,-401,-12,-9,-8,-59,-25,-1,-18,-28,-17,-613,-44,-22,-90,-3,-78,-20,0,-39,-7,-14,-9,6,-267,-1,6,-11,5,-5,-4,-3,4,0,-16,-114,10,5,11,-46,-9,-60,4,-16,13,-2,-38,7,6,-14,-19,-416,-25,-2,-1,5,7,-5,1,19,2,-12,9,-4,-444,-18,-8,3,-427,-20,-10,-5,-21,-8,23,4,-4,-24,18,-9,-10,-43,-26,9,2,-10,-7,-1,-22,-20,-81,-8,8},
{44,51,-2,-21,-30,-5,-10,11,8,1,-2,-11,16,24,-3,-62,-10,-10,6,1,6,4,2,0,-7,-42,-5,-6,47,-107,4,-14,-24,-10,-5,1,18,5,-11,-6,-27,0,19,-22,0,-47,-31,0,2,-6,-32,-12,-48,-36,-18,9,-12,-10,-11,-25,-37,-14,-60,10,-49,-7,2,14,-25,-89,-110,4,-53,4,51,-15,5,35,18,-99,-5,-30,0,6,-45,-44,3,4,-43,19,-38,193,41,4,-15,33,-3,0,24,-20,6,15,0,-185,-7,3,0,-4,-86,-10,7,1,-36,-16,-4,-111,-19,26,-11,-12,-5,-25,-1,20,14,-9,-22,2,-26,1,2,-30,-1,-47,-5,-17,16,5,0,0,1,52,-12,-12,-16,-22,-20,-13,21,-6,-22,15,6,-8,-12,-6,-5,-13,-63,-17,14,8,-31,1,18,6,-26,13,-15,-12,-2,-27,-18,3,2,-13,-42,24,5,-23,-24,21,5,2,-9,-25,-17,5,-2,27,0,22,-12,8,0,-29,22,-48,1,39},
{20,33,0,-36,-77,21,-12,-1,-6,14,10,11,18,28,2,-40,1,-14,30,4,-5,3,-4,12,2,-37,-8,0,59,-46,4,1,-23,1,6,10,15,14,19,4,-37,-1,30,-33,-14,-62,-16,-1,-7,21,-87,-11,-23,-5,-12,20,-16,-3,-32,-34,-40,-47,-81,39,-18,-44,6,24,-24,-64,-75,4,-9,-6,-21,-17,-103,58,19,-120,-8,-43,29,13,-6,-43,10,-3,-33,7,-14,259,54,4,35,42,-7,-9,11,-56,26,-16,-13,-274,-8,-3,-8,-1,-38,-16,24,-16,-27,9,-5,-57,-23,69,5,6,-35,-19,-12,24,-15,-8,11,-31,4,7,-8,4,-3,-16,9,-8,16,5,-1,4,-8,52,-51,-28,0,-77,14,-3,22,-13,-17,0,-3,-9,-21,-3,-10,0,-108,0,16,3,-15,-2,24,-2,-48,18,7,8,-7,-43,-2,4,-3,-27,-49,27,0,-39,-22,49,0,22,12,-59,-16,12,-31,23,4,-3,-3,8,5,-32,13,2,-4,10},
{-43,22,7,-25,-75,25,0,-24,-6,1,8,-1,34,10,13,-29,-3,-10,-14,7,-7,-1,-10,17,23,-29,-5,0,47,-34,-9,40,-17,6,16,22,13,-2,30,-47,-22,-8,11,-27,-17,-44,-18,5,-1,7,-49,0,-8,13,-33,33,-13,-4,-21,-35,-19,-32,-48,46,-14,-33,-12,21,-8,-34,-78,13,5,-4,-39,15,-44,43,14,-98,-3,-50,18,7,19,-33,23,-5,-17,-29,-17,187,64,3,63,36,-1,-5,21,-45,25,-17,-8,-220,-3,2,-5,-12,-73,-21,22,-10,-22,21,7,-40,-6,14,-5,1,-13,-21,11,43,-31,-8,25,-28,-12,9,-3,25,7,-21,-4,4,14,0,6,3,5,61,-64,-39,-13,-13,-7,3,21,-13,-6,-12,-7,-5,-28,10,0,-4,-133,-6,21,-1,-4,8,40,0,-34,29,23,-42,-12,-62,-9,1,6,-30,-42,38,7,-51,-25,46,-11,39,7,-55,-46,10,-39,44,1,-14,-4,17,-4,-31,21,14,-5,-13},
{-78,2,-4,-3,-52,-24,-13,-23,-20,6,-4,-16,52,-23,35,-20,-1,-3,-27,-4,7,1,-9,19,27,-18,-31,-3,49,-19,-8,28,-19,0,33,44,11,15,8,-58,-14,2,0,-15,-23,-29,-29,5,10,3,-45,-19,-10,10,-44,34,-5,5,-26,-54,0,-55,17,36,-5,-1,-1,-2,11,-35,-78,1,13,-4,-36,25,17,-6,5,-73,8,-35,-12,24,45,-21,18,-1,3,-33,-9,138,76,-7,17,28,-9,-15,33,-41,-5,-22,-8,-96,6,-3,5,-38,-107,-9,18,0,-23,28,-5,-7,-22,-37,-8,0,2,-15,25,8,-48,-8,0,-28,-10,8,-6,33,4,-15,14,21,34,-8,-8,2,-4,26,-58,-42,-9,-28,16,11,9,-7,-12,1,6,0,-45,2,4,8,-87,-20,38,3,15,3,45,0,-27,10,12,-43,6,-56,-6,-8,-8,-15,-23,37,-7,-45,-32,29,-7,11,-4,-42,-56,24,-48,59,-4,-25,0,21,-6,-31,32,18,-1,2},
{0,-24,-4,16,-32,-38,-1,-21,9,-20,6,-7,47,-9,28,-7,6,12,-10,2,1,0,-2,48,17,-9,-30,2,28,-7,-4,-46,-22,9,18,49,37,14,-14,-47,-9,5,-6,1,-10,5,-68,0,0,-2,-32,-34,-2,29,-19,36,-19,7,-30,-39,-40,-35,-37,5,3,0,-1,-45,39,-29,-59,6,36,11,-43,7,11,-67,-18,-6,-5,-17,-35,39,57,-3,43,2,6,-3,-8,35,48,4,-32,1,-14,-25,10,-9,-9,-25,4,34,0,-2,0,-31,-121,21,-22,6,-12,16,-3,25,-32,46,-2,-2,10,-17,52,-57,-23,3,-36,-36,12,6,-5,10,0,12,39,0,63,3,-6,1,1,-41,-43,-39,0,-17,4,9,19,0,-22,30,-5,-12,-34,7,-4,14,-18,-1,1,6,41,-8,5,0,-12,3,13,-4,25,-78,12,-7,9,-11,-16,-4,-3,-44,-4,30,2,1,-11,-2,-4,47,0,44,-8,-8,-1,37,1,-10,22,-31,1,12},
{12,-6,2,-11,-5,-23,10,37,37,-33,1,5,45,-8,13,2,10,-4,-8,5,-6,6,-1,-15,21,-35,-34,-8,0,12,-4,-78,12,15,-11,8,0,6,-4,-17,-15,-3,-10,3,17,40,-17,0,-2,5,12,-18,27,20,0,31,-33,4,-8,-56,-22,-27,-44,-2,23,9,-11,-13,64,2,-33,26,8,3,-30,-10,7,-42,-35,-8,4,10,-19,86,66,3,74,6,11,10,3,-105,33,11,15,1,-9,-25,-53,-24,-44,-24,16,-31,4,-2,8,49,-54,38,-44,3,-18,-40,7,8,28,51,14,3,24,-25,52,-63,-24,2,-40,-25,27,7,-5,-6,7,13,78,-5,61,5,-7,-1,2,-25,-29,-1,-18,-10,12,8,32,-33,2,16,-2,-5,-3,-4,-11,25,-58,11,-6,5,41,0,-54,7,-10,-3,-4,-20,58,-81,8,7,0,-10,4,-22,5,-12,36,4,0,-38,-8,9,43,-44,22,17,14,17,1,52,3,-7,17,-23,8,6},
{28,-1,-3,-13,16,-21,-13,16,32,-4,0,-23,40,-3,-15,-24,7,-3,20,7,0,1,-2,-9,31,-79,7,0,-25,-49,3,-47,43,13,22,12,18,-8,-15,15,-21,2,-54,-18,15,34,6,-4,4,24,11,-7,-1,46,5,21,-33,0,-12,-25,-6,-38,17,-40,-4,-4,-6,-9,36,2,10,25,-20,5,26,-12,9,-14,-40,12,-2,43,-1,59,56,33,20,-9,-1,7,-5,-196,0,2,11,-18,6,-24,-88,-14,-62,-16,-11,-28,-2,-1,38,80,8,5,25,6,39,8,1,4,109,-34,8,4,-4,-18,55,-89,6,3,-6,5,59,-2,-2,-13,4,-14,-14,-10,-27,2,-4,-2,1,-69,4,7,-19,14,8,0,39,-4,-46,-15,2,-7,-10,1,37,33,8,-6,-6,-3,42,-2,-25,-8,-17,-11,-14,14,19,-13,-39,-2,-1,16,37,-10,5,-5,2,-5,-3,-1,-52,8,57,-43,20,32,45,70,3,-13,0,-19,5,0,1,0},
{36,-12,-3,3,34,-2,0,-30,28,13,0,-58,31,-16,-10,1,3,-20,0,-5,4,-3,5,25,-4,-67,43,-9,-4,0,-3,-12,37,-51,43,-39,-9,-11,-19,15,-37,0,-52,-7,28,13,62,4,0,-14,30,24,2,3,0,17,-4,2,-29,-5,-68,10,29,-10,7,16,12,35,-8,24,18,4,0,6,18,2,-2,-37,17,39,6,52,1,48,40,9,-38,1,-9,11,-6,-155,-109,-7,-79,-26,-2,16,-107,2,-13,-34,22,-11,4,-2,31,35,16,40,72,4,30,-1,5,-18,65,-6,0,4,22,4,37,-19,-31,8,60,18,11,-3,0,-37,9,-29,-17,-7,-43,-2,5,-2,-8,-84,-10,0,9,-5,0,10,51,16,-16,-4,6,-5,-8,-4,11,-40,14,-26,-5,1,15,1,25,-3,-45,-13,-8,36,-10,45,3,5,-6,-5,0,0,8,28,11,-23,-5,3,-32,5,91,-61,25,30,-12,-19,-4,7,1,12,-37,6,0,-33},
{22,0,2,-23,-2,-13,-14,-74,35,25,-10,-10,34,-17,-27,18,5,-19,-17,0,-7,1,8,40,9,0,32,2,16,-33,-7,12,-7,-45,40,-62,-53,2,11,11,-64,0,7,1,26,-25,23,6,7,6,10,72,5,-32,-22,11,13,6,-4,10,-9,-48,12,-12,-11,21,28,69,-23,-23,-11,32,-12,-3,21,-30,-8,0,41,75,1,28,0,20,13,3,-43,-10,-23,-28,-26,-217,-95,0,-69,-53,9,11,-63,30,26,-48,19,39,4,-5,14,4,-13,42,81,-6,21,-16,-5,-83,59,31,55,17,2,-7,48,16,-10,-3,29,17,17,9,-6,-74,-7,-31,26,-19,1,-4,-4,0,-6,-58,7,-21,37,-11,-50,0,38,15,0,-4,-10,2,4,-4,15,-12,30,10,-1,1,20,5,22,-3,-67,-55,-25,41,-10,21,26,1,-2,-36,-61,6,3,-33,-4,-10,-10,17,4,-13,65,-65,48,20,-80,-92,1,-1,0,51,-65,0,-1,-87},
{19,22,-7,-60,-22,-24,3,-87,27,14,3,35,18,3,-35,41,3,3,-46,-6,3,-10,-6,20,10,8,-14,5,23,-68,6,2,23,-11,42,-51,-76,-14,-35,-2,-31,0,6,1,25,10,-10,0,-2,8,-5,53,-18,-33,-74,-24,14,-8,1,0,-20,-96,-27,-25,-81,15,38,47,-37,-39,-26,46,-32,2,38,-40,0,13,29,58,6,42,10,-4,-38,-6,-7,-11,-28,-47,-9,-66,-76,0,7,-54,3,-13,-35,46,40,-36,16,28,7,0,-17,0,-8,25,50,0,12,-7,5,-99,14,63,33,12,-1,-42,-1,0,-4,5,-1,1,7,0,5,-24,-2,-35,23,-36,14,0,-4,-4,-5,-11,15,0,28,1,-24,-14,25,27,-12,-56,7,14,-24,0,-9,14,23,0,-17,-5,28,-2,29,3,-103,2,-21,12,-13,24,76,-7,0,16,-41,-4,-5,-11,-21,25,-2,76,10,-6,43,-29,27,4,-132,-94,-4,-11,2,42,-45,21,-10,5},
{14,6,6,-59,-7,-26,-26,-86,12,10,5,21,0,0,-16,34,2,-34,-36,-4,-2,-7,-5,15,17,19,6,-4,36,-65,1,9,52,-2,55,-32,-57,-7,-51,-4,-25,6,-7,-7,29,22,-22,4,-3,23,3,52,-27,13,-18,-12,-34,3,-1,-15,-46,-70,-43,-2,-85,4,26,23,-31,7,-7,34,-58,-12,-1,-12,-15,10,29,0,6,1,2,-18,-70,-10,-9,-1,-14,-85,3,-37,-30,0,13,-9,-4,17,-71,27,61,-20,1,15,2,-12,-23,-16,-7,19,-12,0,17,0,-3,-73,68,58,-12,10,5,-52,-33,-29,42,-1,-9,3,36,0,1,0,-7,-85,34,-35,20,2,-1,3,-6,15,0,-8,-59,7,0,-7,20,16,-11,-67,1,6,-19,-16,-26,40,-5,7,-14,3,26,-1,50,6,-178,8,-21,16,-5,18,32,2,-8,11,-2,-22,-7,19,-4,44,-3,44,10,-5,15,-52,-9,-10,-162,-66,-6,6,-1,-2,-29,6,-4,47},
{7,-42,0,-37,-19,-10,-20,-63,12,3,-2,4,-24,-18,-10,19,-6,-37,-21,0,4,0,-11,-1,18,17,17,-6,1,-6,2,-9,65,-5,37,4,20,-15,-44,-12,-1,2,-3,-16,10,7,-28,-8,3,21,-5,23,-3,54,48,0,-34,3,-23,-5,0,-4,-25,-8,-71,-5,24,6,-23,-24,-21,6,-29,2,-105,-4,-25,-16,4,-62,-4,-4,4,-40,-102,5,-10,-6,3,-74,0,-11,-5,-2,11,18,-10,-61,-104,2,47,-17,-16,-27,0,-1,-32,-22,-20,-17,-65,6,0,-6,4,2,8,27,-26,-18,-1,-26,-26,-44,9,3,-8,-4,12,3,2,20,5,-46,24,-22,28,2,-10,-3,5,-16,-11,-3,-115,-6,12,-10,2,-5,-12,-12,1,1,-18,-11,-18,30,-2,0,-20,5,10,-3,48,8,-44,8,11,12,-2,-4,27,-4,-3,5,32,-36,-6,11,-1,42,-1,34,7,-2,22,-42,-9,-4,-21,-50,0,-3,1,5,-27,1,-6,31},
{-113,-58,6,-14,8,6,0,-16,-27,-45,-1,0,-20,-18,-7,2,-13,10,4,-1,-4,-7,0,-8,-4,-23,-26,7,-35,-13,0,-74,-3,3,-4,-5,8,-29,-15,5,1,7,3,-69,-17,-45,-13,-1,3,-4,-19,-3,13,4,16,11,18,-6,-22,-21,47,7,-14,-27,-3,-52,-14,-46,-20,-12,-18,-13,7,-9,-31,24,9,-5,2,-2,6,-5,-5,7,-44,-20,-1,-7,-15,1,7,-518,-1,-2,4,-12,-22,4,2,1,-24,-26,-45,17,3,-1,-16,-1,-124,-79,-20,-14,-51,-14,-5,-7,-13,4,-10,-64,-13,17,3,-10,14,2,-40,6,-3,-8,-8,-8,3,-30,4,2,7,-5,-3,-5,4,-2,6,11,-3,-6,-11,-18,-20,10,0,-5,5,-21,-2,-16,4,-1,14,-16,-42,0,-30,-6,-5,-2,-3,14,3,-21,-6,-23,-12,4,0,8,4,-22,0,-14,-8,-21,2,0,-30,-11,-41,-7,-72,1,-7,-8,-12,-13,-8,-20,-10,-1,0,-28},
{-11,-11,7,-3,-6,-5,-6,-67,-6,-14,-1,6,-33,-6,-527,-49,-4,-7,-7,3,-7,3,1,-33,-8,-115,-1,-1,-8,0,-9,-15,-7,0,-16,-77,-69,-202,-9,-7,-6,-8,0,-39,0,-3,-10,0,-3,-2,-7,-11,-84,-9,-10,-5,-7,0,-18,-12,-3,-11,-15,-49,-66,-42,-16,-6,0,-10,-17,-18,-2,0,-2,-2,-18,-17,-3,-11,0,-76,-12,-21,-48,0,-6,-5,1,-14,-33,-15,-13,-6,-3,-10,-16,-10,0,-4,3,-19,-25,-11,3,4,-4,-7,-268,-8,-8,-2,-7,-5,-3,-121,3,0,-12,-43,0,-11,-8,-6,-10,7,-17,-14,-10,-4,-1,-63,3,-8,-2,-10,-1,6,5,2,-3,2,-8,-6,-16,-14,-15,-2,-22,-15,-5,-12,-5,-165,0,6,-3,-13,-15,-14,-7,6,-16,4,-89,6,-5,-4,-14,-11,-42,-14,-11,-9,6,-3,-7,-11,3,-9,-4,-35,1,-7,-121,1,0,-19,-20,-18,-12,-41,-11,-9,-2,-5,-7,-14,-2,-6},
{-5,24,6,-30,9,-6,-13,-17,-32,6,6,-31,23,18,1,-12,-10,-11,13,-6,4,-1,-1,2,-11,-60,-30,-6,24,-48,-3,-15,-78,-11,-8,8,15,0,-16,-16,-16,6,15,-36,-14,-28,-28,-7,-6,-24,-28,-21,-57,-66,-11,-6,-5,1,26,-140,17,10,-16,13,-16,-2,-4,-5,-19,-32,-46,-11,-29,3,42,-27,-16,27,4,-29,-8,-18,-3,14,27,-15,1,6,-27,-9,-13,118,31,2,-5,-547,-17,-4,19,-10,-20,-13,-9,-111,-9,-8,-6,-66,-132,-24,-16,0,-1,-21,-4,-69,-10,9,-77,-41,1,-39,-2,23,-8,-6,-6,20,-57,0,0,-23,5,-90,-5,20,8,-3,0,-5,-7,31,2,11,-25,-8,-49,-22,7,-1,-16,4,0,-29,-7,-11,-2,-7,-29,-14,24,3,-17,-7,3,2,2,11,4,-31,-15,-17,-24,-9,5,-37,-13,12,2,-26,-175,9,-3,4,-28,-20,-6,22,-25,29,8,-3,-22,0,7,-29,14,-45,1,23},
{-8,26,-2,-31,-11,4,-5,-30,-58,3,-7,-6,42,16,6,-11,-19,-7,-6,-5,4,3,-3,3,-17,-62,-11,-8,23,-21,4,27,-44,-17,10,28,10,-1,23,-24,-19,0,27,-42,-14,-27,-41,-5,3,-15,-67,-6,-94,-60,-57,-16,9,7,-5,6,8,30,-33,30,-15,0,-23,18,-9,-42,-44,-3,-3,-6,-5,-36,-32,40,1,-73,-1,-24,10,28,45,-7,8,-4,-37,-10,-16,200,44,3,-14,50,3,8,42,-39,14,-12,2,-53,-2,-8,-22,-41,-103,-42,3,-1,-16,-1,3,-77,5,94,-62,-22,-17,-40,0,35,0,-8,10,2,-54,1,-7,6,-5,-101,0,58,-11,0,-2,4,0,42,0,-21,-34,-44,3,-1,41,-15,-24,-24,2,-15,0,-8,31,-20,-50,1,13,5,-10,0,21,1,5,-4,-8,-32,-60,-18,-11,1,-1,-19,-18,26,4,-42,-73,11,-8,24,-25,-37,-22,36,-31,38,19,-16,-4,0,-7,-38,-11,-41,6,16},
{0,16,6,-11,-48,2,-5,-42,-50,0,5,-14,46,9,19,-6,-11,-10,-5,-1,-6,-8,0,0,-1,-30,-5,-5,29,-34,-2,40,-24,-7,18,21,0,1,34,-37,-17,-9,30,-44,-18,-29,-43,0,-5,0,-53,-20,-98,-41,-60,-4,-3,0,-25,7,0,16,-60,18,-15,-12,-2,20,-2,-33,-33,1,34,-12,-9,17,5,9,-5,-85,-3,-25,2,33,42,14,21,0,-28,-4,-16,201,43,-12,44,16,-9,0,34,-57,14,-6,0,-124,-3,-5,-19,-19,-101,-19,1,-6,-24,33,-1,-74,9,103,-4,6,7,-35,3,31,-2,-3,0,-37,1,-6,-6,13,-10,-34,5,96,-2,5,0,-4,6,40,-16,-18,-29,-28,38,2,42,-14,-8,-17,-2,-35,4,-10,23,-15,-103,-2,7,1,0,-4,29,3,4,-8,5,-18,-58,-15,-6,-7,-2,4,-14,9,1,-38,-49,-21,5,29,-18,-45,-29,12,-43,33,21,4,-9,7,8,-29,6,-3,1,4},
{35,15,-3,11,-46,-14,-11,-38,-10,-7,1,-26,55,-7,29,-11,-3,-8,-20,8,1,-6,-7,11,-8,-33,-7,3,31,-39,6,-8,-29,-1,28,23,-19,19,19,-38,-20,-3,13,-9,-6,-9,-94,0,-3,8,-12,-5,-98,-29,-76,4,-19,-1,-23,5,-12,22,-44,23,7,0,5,5,5,-21,-36,21,42,-4,-61,27,18,-19,0,-69,8,-28,-17,45,44,18,36,2,-24,-7,7,168,45,2,34,5,4,1,31,-32,0,-1,20,38,1,0,-23,-52,-100,14,-7,-6,-11,47,-10,-52,-23,77,14,20,26,-31,2,-1,-4,-6,-65,-33,34,-6,-9,14,-8,14,20,93,8,6,1,-5,0,12,-21,-35,2,-23,57,-2,39,5,19,17,4,-42,-22,-1,21,-5,-57,1,2,-4,5,8,20,0,-31,-23,-11,-32,-11,-23,1,3,-2,27,-17,8,0,-39,-49,-79,-4,18,-39,-23,-19,20,-12,34,-1,-1,2,23,8,-21,34,2,0,0},
{35,6,1,35,-1,-16,-6,1,33,-13,1,2,37,-44,32,-8,8,7,-10,-8,0,-5,10,26,-15,-37,-23,4,21,-35,-8,-77,-29,-4,-6,19,0,13,14,-18,-4,-9,-8,2,8,30,-53,5,-4,-5,0,-18,-76,-24,-54,0,-48,-8,5,-12,-20,-32,-102,-23,6,34,11,-1,24,0,-27,35,40,-5,-35,16,13,-29,-31,-33,-4,-17,-43,47,34,6,80,5,-9,12,13,1,33,-7,-27,7,0,-4,19,1,-14,-9,49,-36,4,4,-10,-9,-81,48,-39,-6,3,24,-12,-33,-11,54,28,30,44,-18,6,-68,-2,-7,-47,-23,36,3,5,9,-3,27,57,-22,53,-8,1,4,1,-51,19,-36,9,-4,30,0,45,12,16,35,6,-36,15,-7,-62,19,-73,20,28,-3,27,0,-40,-2,-13,-53,-19,3,35,-63,21,6,1,45,-12,-9,3,-26,15,-115,-4,32,-36,-7,-22,19,-2,35,-5,-8,6,64,-8,-23,29,-11,-8,31},
{18,-8,9,15,-20,-15,-8,-22,27,-24,1,33,28,-14,14,-16,-4,12,-5,-1,8,4,-2,-33,6,-44,5,-3,-41,-40,-4,-17,-6,10,-16,-8,31,16,20,7,-2,-7,-16,9,12,45,25,-7,7,3,6,-23,-51,-17,-22,11,-44,-5,-45,-38,-16,23,-85,-18,23,36,10,30,39,3,-7,50,18,0,-2,-16,18,-14,-50,0,3,7,-17,63,35,0,44,-3,-8,17,17,-105,15,1,-87,-1,-3,3,-46,-7,-9,-32,49,-36,-8,8,-22,25,-52,52,-41,-1,-46,-23,-10,-29,23,34,42,36,27,-11,0,-77,-6,-5,-10,-2,30,-4,-8,7,-7,19,78,-25,46,-7,-8,7,6,-70,23,-4,-12,-17,8,2,58,11,6,1,-4,-3,5,0,-40,29,-67,44,32,-2,15,-5,-62,0,25,-40,-27,2,64,-44,4,0,2,46,-14,-9,5,-16,40,-129,-4,42,-27,6,-33,-104,17,35,16,5,1,26,2,-15,29,-1,0,51},
{3,5,-3,-5,2,6,-16,-52,21,-32,-2,11,21,-27,6,-15,-5,14,-18,-2,-8,-7,0,-21,20,-113,38,-4,-32,-99,4,-7,-4,31,12,-50,-1,5,-5,30,5,-6,-24,-7,15,48,30,-8,6,22,25,-15,-51,-27,-16,5,-4,0,-43,-1,17,39,-2,-5,15,28,21,5,2,3,17,55,-3,-8,28,-9,16,4,-16,13,0,28,16,45,22,-15,-6,5,-2,20,16,-152,-23,-10,102,-18,-7,23,-110,-13,-28,-21,13,-32,0,-4,6,44,18,25,-8,8,5,22,-12,-25,65,-25,-26,11,4,-15,-7,-14,-15,-9,-24,-1,32,-4,5,0,0,27,0,-29,-26,-3,-4,-2,-4,-81,24,15,-43,3,9,-5,55,-9,0,-22,3,13,-32,5,-13,18,2,13,0,1,23,3,-6,-3,-5,-18,-29,22,56,60,-24,0,-1,92,-34,-18,-4,-6,8,-87,-6,68,-91,9,3,-86,11,41,22,19,0,-32,2,-17,3,1,0,44},
{18,-15,6,14,17,1,-13,-87,4,23,-1,8,29,-24,-14,3,-7,-8,2,3,-4,-4,3,13,-10,-84,42,0,-2,-58,-9,8,0,-34,57,-81,-31,-12,-17,28,1,2,-19,-2,4,37,19,-2,-9,9,20,-1,-27,-2,-15,10,6,5,-9,-14,-59,80,-10,-25,13,23,25,38,-6,11,12,22,3,4,23,2,5,-11,17,30,6,22,-14,44,16,-40,-51,-8,11,26,15,-168,-113,0,-28,-19,-6,48,-112,0,-37,-14,13,1,-9,-7,21,18,7,10,10,5,4,5,-8,-22,88,-1,-41,20,14,-5,17,60,-14,-6,45,0,-1,7,7,-39,-5,-14,0,-3,-61,2,-7,-2,-6,-77,21,6,-25,-10,2,0,56,8,22,-35,3,0,11,-8,1,-40,16,4,-6,1,2,5,33,-2,-33,-16,-40,33,5,45,-27,3,-6,5,-39,-5,-6,18,1,-84,-8,29,-34,2,35,-72,6,37,17,-28,15,-23,0,11,-20,14,0,21},
{6,8,-7,-5,5,-3,-33,-112,3,17,-8,-3,22,0,-30,14,-8,1,-12,-3,6,-2,-6,6,5,-3,8,3,4,-37,5,12,10,-55,57,-101,-87,-9,3,19,-31,2,-1,5,12,-10,6,-4,-2,11,13,17,-6,-26,-11,9,5,-8,10,-6,-19,-32,8,-50,16,16,33,44,-7,-4,-10,33,-2,4,59,-8,-10,4,35,17,-8,14,-21,6,-13,-28,-43,1,7,-23,-18,-178,-99,-13,-28,-44,8,47,-15,11,57,-15,2,17,-3,8,3,5,-7,28,5,-6,0,1,-6,-57,74,32,38,19,1,-6,8,27,2,1,10,21,4,6,-9,-104,-7,-21,42,5,-5,7,0,4,5,-28,10,-23,11,-10,-22,-14,27,19,0,-24,-5,4,6,-20,1,-46,8,9,-1,-4,18,6,44,-5,-40,-27,-57,14,-22,16,-26,7,8,-18,-57,2,3,-5,2,-33,0,56,13,-6,4,-19,21,30,-43,-106,6,-14,-5,33,-35,0,-2,-29},
{3,0,5,-28,-25,-24,-16,-105,11,6,-6,21,-4,4,-44,46,-3,7,-53,1,2,-9,-8,-15,11,2,-10,6,19,-57,-2,21,27,-13,46,-90,-94,-20,-25,20,-33,0,-4,-4,27,24,1,-10,5,12,-19,24,-15,-12,-51,-14,22,-2,8,-19,8,-3,-24,-52,-11,6,17,23,-8,-50,0,19,3,3,50,-40,-14,12,31,18,3,-1,11,-20,-65,-52,0,-4,-23,-35,-8,-55,-46,-13,12,-36,9,31,-11,6,22,-14,4,2,0,-7,-6,-20,6,10,-4,-9,7,12,2,-90,37,29,4,1,-23,-19,11,16,4,-10,-6,0,36,4,-5,-32,2,-26,34,-27,16,0,6,-7,6,-11,3,-12,9,0,23,-19,33,13,0,-65,4,9,-14,-3,-21,5,6,-8,-23,6,22,-8,34,-7,-110,-8,-13,15,-13,13,-6,1,-8,12,-44,4,0,1,-18,24,6,58,2,7,9,-29,12,4,-89,-50,-1,-20,-13,31,2,4,3,-14},
{3,-25,-4,-50,-25,-31,-18,-81,0,8,0,8,-4,-8,-21,32,-6,-6,-33,-6,-5,0,-2,-5,18,10,-9,2,20,-42,-4,6,27,16,36,-47,-52,-30,-41,0,-2,0,-12,-13,24,20,-10,-5,-8,36,-26,30,-34,49,-32,-21,4,-3,7,-23,-6,40,-38,-37,-46,-3,6,-3,-17,-50,-3,25,-17,-4,-22,-19,-15,-5,13,-14,6,-18,3,-36,-81,-53,11,-8,-16,-39,5,-29,9,0,14,15,-9,25,-41,4,19,-12,-14,-6,2,2,-24,-36,5,-16,-70,-4,1,12,-5,-61,16,18,11,-7,-13,-40,-15,-8,0,-5,-11,-3,24,-4,4,-1,0,-78,34,-23,28,8,-7,3,3,-8,0,10,-35,3,5,-21,19,0,11,-28,-8,5,-34,-17,-28,20,-5,-14,-27,-2,35,0,37,0,-79,6,2,8,-14,-5,0,5,-2,25,-2,-18,4,-9,-13,32,0,0,6,6,10,-21,1,-2,-34,-27,-1,-8,-14,-2,13,10,1,9},
{0,-18,-8,-31,-35,-10,-8,-58,-2,3,-1,-31,-13,-33,-54,21,-3,-31,-17,8,6,0,0,-29,37,14,-13,-5,16,-24,4,16,35,15,28,-39,-63,-40,-29,-7,-5,-1,-12,-25,13,14,-31,-8,-6,11,-14,22,-41,31,-11,0,-22,0,-21,-13,4,8,-32,-97,-84,-17,22,-21,-12,-23,-15,26,-50,-8,-27,-2,-31,-3,7,-35,8,7,9,-64,-106,-37,15,3,1,-39,18,-13,-1,-5,8,12,-11,-52,7,3,3,-19,-23,-70,3,-4,-57,-12,15,-77,-59,1,-1,0,4,-9,19,19,-21,-19,-23,-25,-20,56,13,3,-24,2,-9,6,5,2,0,-53,47,-10,30,-6,7,0,2,-29,-20,8,-32,9,-2,-6,14,11,29,-4,0,-14,-28,-4,-20,5,-3,-21,-12,6,33,-4,-11,0,-34,20,13,12,-20,-8,10,1,8,36,14,-29,0,-4,2,19,-5,23,-3,11,11,3,-16,-12,0,-1,-24,-13,-12,-19,-20,3,-4,0},
{-26,-10,-7,-3,-1,-5,-1,-278,-15,-112,6,-304,-20,-7,-79,8,-14,-20,3,5,-1,-9,-1,-17,15,-18,-44,-8,4,10,-9,-1,13,8,-24,-60,-463,-53,-3,-1,-2,2,-1,-58,7,-14,-2,-6,-6,-20,4,-32,-1060,1,1,1,-8,-5,-13,-101,-118,-71,-6,-2,-156,-30,7,-21,-27,1,-18,-38,-4,1,0,-2,-1,0,5,0,-6,2,9,-36,-558,-343,-2,-3,7,-96,-7,-38,-6,-7,-398,-43,-16,21,-19,-45,-250,-11,-40,-109,0,-9,-11,-7,-30,-33,3,4,-31,-7,4,-34,9,-646,-415,-32,-16,1,-11,-1,-14,5,-18,-5,-84,0,-2,-18,-7,28,10,0,3,-6,6,0,5,-20,-8,-1,7,1,5,-11,-8,-21,14,13,1,-41,5,-1,0,-24,-24,-34,4,8,3,7,-108,6,6,-2,10,4,0,-17,7,-3,-1,15,-31,-2,0,3,-3,-67,0,16,-25,1,-48,-944,-48,-12,26,6,-23,1,-3,8,-24,-19,-1,-308},
{-10,-1,8,-3,-5,-7,-1,-62,-7,-5,-7,3,-19,-10,-523,-41,-6,-7,-5,-4,-3,2,-5,-32,-8,-117,-6,-8,-5,-12,0,-13,-2,-11,-25,-66,-69,-171,-4,0,-11,-9,-1,-49,-12,-15,0,4,-10,-3,-8,-11,-85,-10,-13,-8,-8,5,-15,0,-8,-9,-6,-57,-63,-39,-18,-12,-2,0,-20,-21,-3,0,-11,-4,-30,-1,-5,-12,-4,-81,-11,-17,-65,-6,-8,0,2,-7,-48,-6,-17,0,-13,-8,-15,-19,-7,-15,-6,-17,-26,-7,-7,-1,-10,-6,-241,1,-5,-10,-8,-13,-6,-112,-1,-14,-7,-45,-13,-12,-10,-6,-6,-7,-5,-3,-11,2,0,-65,3,0,-19,-7,-8,-8,-4,-9,3,-5,-4,-4,0,1,0,-4,-29,-22,-11,-12,-5,-158,-1,5,-14,-12,0,-28,-12,1,-8,5,-77,0,-11,0,0,-13,-27,-26,-1,0,8,-7,-13,1,-3,-17,-7,-28,-10,-10,-115,-3,0,-25,-18,-22,-16,-29,-12,-10,5,-16,-20,-24,0,-7},
{-143,0,-2,-11,-9,-7,-8,-87,-47,16,-3,-124,-11,-1,-45,-2,7,-3,-3,-8,-6,3,-3,-4,-11,-102,-1,-2,-7,-9,0,15,-187,-7,-5,-285,3,-56,0,0,0,2,-4,-57,3,0,20,6,6,-4,-37,-9,-31,-8,-13,-12,0,-8,-32,-13,-12,6,20,-8,-11,-19,-36,-6,-12,-3,-11,0,-12,3,-10,-157,-36,-2,-2,-4,-6,-21,-2,-18,-30,-310,-6,8,-21,-2,-11,1,-3,-9,-12,-12,-9,16,-541,-37,-30,-30,-10,-16,-4,-11,-14,-176,-1095,3,9,-7,-6,2,-9,-30,5,-12,-84,-25,8,-20,-12,-83,1,-9,29,2,-28,0,5,-39,-7,-223,-4,-62,1,0,-7,6,-7,13,-4,-5,-25,-7,-17,-18,-20,-32,-6,-11,-2,-184,-4,-10,12,-4,-1,-17,-1,8,0,-4,-16,0,-7,0,-51,-16,-345,-18,-4,8,-8,-18,6,-4,0,-13,-413,-75,-1,1,-492,-27,5,-2,-14,-16,-2,-174,-26,-1,-10,-2,-12,-50,0,-15},
{-22,-22,2,-22,-176,-28,-7,-62,-53,-9,1,13,-30,-43,7,5,-5,-6,-25,0,-3,-1,1,11,-31,-118,-5,3,1,6,-6,41,-45,-8,1,0,-35,-5,-26,-43,-33,0,-2,-28,-19,-16,-38,5,3,-17,-55,-29,-112,10,-14,-31,-15,-6,8,-366,-22,31,18,7,-3,-20,-96,-27,-8,3,-4,-14,-4,4,-11,-41,-73,-16,-5,-9,0,-28,-15,-25,-35,-11,-5,-6,-27,-18,-19,56,19,-2,4,-5,-4,20,-25,-79,44,-50,-11,-40,-1,0,0,-57,-377,-15,18,7,31,28,-7,0,34,-5,7,-36,-12,-5,-27,11,-17,0,23,-28,0,-2,-3,-29,-4,-246,-7,23,-7,-6,7,-5,1,-25,-29,-31,-98,-31,-9,-17,-22,-23,-25,-90,0,-135,-29,-8,28,0,-37,-3,-10,5,-9,-2,4,0,7,-2,1,0,-199,-404,9,0,1,-131,8,-14,1,-17,-116,-317,0,23,-737,-59,-24,28,2,-34,24,-69,-12,1,-6,0,2,-56,1,41},
{-30,-26,1,-13,-2,-8,-14,-55,-39,4,3,-4,-20,-27,19,3,3,-2,-23,-3,-7,0,-7,15,-28,-54,-1,-3,12,-21,-1,25,-65,-4,7,50,-158,16,-14,-34,-22,0,-2,-2,-16,-31,-102,-1,-2,-8,-24,-28,11,37,-10,-21,-4,-4,-55,-210,-55,15,13,5,-3,-24,-52,-25,-4,-6,-11,0,6,-1,-52,-3,-61,-11,0,-18,3,-19,-24,-21,-23,109,8,5,-25,-19,-6,46,23,-7,-23,-3,-16,7,8,-54,55,-29,-10,-86,7,0,-19,-26,-350,0,19,0,18,36,-6,7,31,17,19,-9,-15,-42,-3,62,-10,2,-31,-38,12,4,2,4,-5,-111,9,17,-1,3,-9,2,0,-32,11,-19,-117,-18,16,-8,-13,-35,-21,-97,3,-185,-27,2,30,1,6,-6,-12,-2,6,7,17,0,4,-11,-16,0,-280,5,16,-3,-5,11,8,-20,-8,-38,-128,-17,-2,20,-84,-36,-26,31,-2,-12,16,-79,1,13,1,-3,-2,-46,-2,22},
{12,-12,0,-11,13,-13,-33,-18,-6,-1,-7,-15,-9,-23,19,2,0,0,-12,5,5,2,-3,13,-10,-116,9,-2,16,-42,7,-52,-51,-6,8,13,-191,11,-10,-4,-3,-8,-9,2,-12,-5,-184,1,-3,0,-29,-14,33,48,-16,-6,-34,5,-28,57,-113,6,0,-20,-2,-19,-73,-18,-3,-4,-2,-4,-6,-2,-92,-22,-24,-10,-10,-18,-5,-10,-8,-1,-19,105,17,-7,-15,-8,15,40,15,-1,-40,54,-4,18,6,-34,34,-11,-13,53,-4,3,-12,-41,-163,19,-3,-6,50,33,-2,5,14,50,22,-19,-6,-12,-14,48,0,-7,-114,-29,16,-6,-7,56,3,-48,26,-12,6,5,-5,0,-5,-34,28,-17,-19,-18,14,-10,5,-35,2,1,0,-159,-23,-7,22,17,48,-6,-10,-1,2,-8,-17,3,-53,-21,-43,-18,-45,-270,22,-5,-5,7,6,-10,-5,-18,-50,-68,7,25,-51,-24,-27,40,-4,-56,9,-101,-9,18,-3,-10,15,-32,6,4},
{4,-3,3,3,20,0,-26,-38,-3,5,-4,36,2,6,6,-20,-24,-1,-9,-7,1,-1,0,7,-8,-54,-21,-6,22,-21,-5,-105,-72,1,-44,-41,-60,2,38,0,8,7,6,9,14,5,-53,0,2,-17,-4,-36,7,-9,-8,-1,-49,-4,73,-2,-6,20,-68,-58,10,-1,-36,8,-1,-4,-1,0,-8,-7,-25,-7,-9,-14,-34,-6,-2,4,-3,29,-27,1,23,-9,-11,-1,3,1,2,-2,-52,21,-10,48,19,5,24,0,3,0,-5,4,-32,5,-41,11,-14,0,25,-3,-7,14,44,25,3,0,4,-4,0,28,-12,1,11,-8,12,0,4,52,-9,-47,32,-34,35,-2,-7,0,1,-75,30,-8,-19,48,7,-12,14,-5,-15,10,-6,-152,35,-14,-33,10,-16,0,10,-4,23,2,-91,7,-67,-7,-14,0,118,-257,25,0,-7,-4,6,-10,-9,-5,6,-106,-10,48,-5,-1,-3,8,0,-16,0,-48,2,33,-3,-11,3,-18,-3,26},
{-7,-13,5,4,22,-7,-8,1,6,-10,-8,16,11,-8,-35,-32,-25,4,9,0,4,5,-12,-29,6,-29,-11,-1,26,-151,-2,-66,-86,-11,-68,-73,25,-19,4,16,-2,0,-9,7,-17,-4,18,-1,-6,15,-14,-12,-3,2,0,-12,-21,7,-18,-7,17,-18,-37,-59,20,1,4,-4,-21,0,-2,8,-5,4,6,0,2,1,-39,-7,0,5,-5,-3,-2,-42,-9,-1,-8,6,21,-41,15,-9,4,-12,-3,45,-14,-6,38,7,0,-21,-1,-2,-2,3,-8,4,-11,8,0,-7,3,14,58,4,0,-7,5,-1,-22,27,0,-6,73,-9,-3,-2,5,-20,3,1,24,-24,38,-2,-1,-8,-4,-71,4,5,-50,31,0,-11,-12,-3,-35,-43,-1,-86,-8,-1,-19,12,-13,-8,-7,4,48,-7,-116,4,29,11,-160,-7,118,-80,10,7,7,-41,0,-8,4,1,-1,-83,2,51,-90,2,-20,-23,6,18,8,-16,-9,15,0,-14,4,4,7,24},
{-15,-1,1,5,4,-3,-6,9,2,-25,4,-7,9,-27,-61,-9,-22,1,-3,2,4,-6,0,-14,7,-82,-14,7,11,-59,6,-15,-74,-6,-49,-79,-8,-59,-19,0,-5,3,-14,0,-15,-1,27,1,7,16,3,-20,-21,-1,-11,-9,20,-1,-37,0,18,-1,-10,-38,16,8,45,-14,-69,-14,0,0,3,-6,23,3,5,-26,2,-6,0,9,-3,-29,-9,-62,-37,-5,-11,0,3,-83,-22,-10,62,-20,5,7,-14,-2,54,15,5,-7,7,-8,-9,-4,27,-9,52,-11,2,59,3,21,71,-20,-16,-11,-5,-9,-7,36,-10,6,68,-2,-9,-2,-1,9,0,17,-64,3,-25,2,3,6,6,-39,13,3,-72,12,-3,-17,-13,-6,-25,-110,4,-8,-24,0,-5,-8,1,-12,-26,0,36,0,-67,6,0,-10,-23,-20,51,44,-16,0,-8,-3,0,5,0,0,-6,-35,1,87,-153,11,-22,-31,-8,9,42,-53,2,-24,-2,-26,-4,2,1,26},
{-6,-35,0,8,0,16,-6,32,-16,4,4,-135,21,-21,-55,-9,-16,-7,-15,3,4,0,3,-41,-27,-37,-5,-10,-40,-7,3,-5,-19,-18,-57,-24,37,-77,-27,-17,-3,-4,-4,10,-8,-3,11,-5,-6,-14,21,-25,-40,1,0,1,14,1,-13,8,-49,13,-3,28,17,7,41,0,-53,0,3,-39,2,5,23,9,3,-15,7,0,-8,14,-21,-44,-14,-14,-6,-5,-12,-8,-6,-110,-88,4,-29,-15,5,55,-23,0,-14,12,0,-3,1,-10,9,-9,25,-50,-5,-8,1,40,3,13,39,-6,-42,-3,-6,7,9,45,-25,-2,-5,8,-27,1,5,-67,-8,-7,-39,14,-16,3,7,-4,4,-94,4,-14,-29,-11,-12,-11,0,0,-42,-109,7,2,1,0,21,-45,1,4,-17,1,1,-5,-44,-1,-67,-24,-19,27,-5,9,-33,1,-6,-24,-11,-4,-9,10,-1,-87,-10,70,-77,-2,-20,-54,-2,6,18,19,-3,33,-2,1,-1,9,4,-18},
{-4,-57,7,-8,-4,8,0,-63,-29,-5,7,-150,-6,-14,-55,6,4,-3,-2,0,-8,-8,-7,-68,-54,2,-13,3,-38,4,-2,18,-25,-50,6,-46,21,-70,-22,-3,-8,-7,-11,2,-4,-13,3,0,3,-1,0,-64,4,25,-7,9,0,5,-5,-8,-19,27,-12,9,12,-8,71,2,-27,-9,-4,-24,2,-5,55,6,-6,-18,16,3,-8,7,-41,-6,-26,-100,-2,-6,-14,-32,-21,-30,-105,5,-16,-6,0,55,-9,0,-115,4,0,9,0,-3,-10,-5,27,-47,6,0,4,76,0,-5,8,0,-25,-11,-6,0,8,13,-20,1,-43,9,-39,2,-5,-128,-1,-26,16,15,16,1,2,-8,-7,-30,0,-24,-34,-14,-4,-10,-4,-1,-79,-38,-2,-9,-7,0,10,-75,1,-1,-1,7,7,0,4,-5,-64,-21,-38,-46,-117,-1,-29,7,-1,-79,-11,-8,-7,-2,-9,-41,5,40,-7,5,-5,-17,-2,-13,15,-6,0,25,1,50,-10,6,-4,-9},
{1,8,6,-4,-2,3,-1,2,-73,-4,-2,-366,-43,-12,-34,31,1,-5,0,0,-4,6,0,-70,-32,0,-1,0,6,0,2,13,27,-44,-6,-85,31,-89,-29,0,-53,-6,-20,-7,-14,-28,5,7,-1,15,-1,-73,-53,31,-3,-23,-3,7,7,-2,-4,0,-34,-29,10,-20,37,-21,-11,-32,-5,4,-9,-9,26,15,-18,-11,31,0,-8,-33,-11,-34,-16,-95,12,-3,-26,-26,-65,6,5,6,5,4,10,11,-34,-8,-378,9,3,9,-4,-3,8,-6,29,-56,-21,-9,-5,51,-2,-78,7,-3,-29,-17,-44,-4,10,-11,-18,-3,-64,-15,42,7,-4,-67,3,0,11,11,1,6,3,-4,6,-18,1,-18,-81,2,22,-7,-57,3,-42,-72,-2,0,-32,-6,-11,0,5,-12,-11,0,0,2,1,8,-71,-56,14,2,-75,-9,-11,-1,2,13,-44,-11,5,-51,-18,-6,1,15,-10,-13,-9,18,2,40,22,27,-5,-18,-3,31,6,20,-8,-50},
{9,-16,5,-40,6,-10,-2,-93,-172,-1,-3,-768,-117,-36,-69,4,5,-34,9,0,-7,-2,2,-68,12,3,6,5,11,-73,-1,34,-15,3,8,-100,-23,-93,-40,-23,35,4,-46,-8,8,-4,-6,0,-2,-14,-73,-14,-90,-1,-6,-14,-31,4,-7,3,-16,16,-44,6,12,-23,-57,10,3,-14,-11,-3,-43,0,-47,-5,-9,-24,1,-2,0,-27,20,-187,-37,-400,9,-5,-25,15,11,20,6,2,2,34,-13,35,-248,-3,-404,0,-6,-7,2,-4,0,-24,22,-79,5,-18,6,23,1,-18,2,0,-9,-22,1,-4,10,-262,-8,-4,-115,-28,-15,3,-9,-14,0,-172,14,9,12,1,1,5,6,-12,-4,0,-46,-6,21,-14,-150,-2,-22,-12,0,-10,-33,-6,-28,8,-10,-12,8,-9,9,1,12,-8,-1,13,43,-29,-809,-20,5,-1,-7,35,1,-58,-5,-11,-52,-43,1,13,-17,15,12,35,6,-7,20,-15,-1,-40,5,-14,1,-12,1,-12},
{8,-11,2,-45,-274,-11,5,-807,-66,7,1,-24,-32,-35,-56,11,-18,-27,-22,-4,-4,1,-3,-9,-17,-1,11,-5,14,-148,0,24,-71,-9,16,-264,-47,-66,-47,-19,-23,2,-19,-13,2,-7,-85,-4,3,-4,-78,5,-171,0,-14,-22,-77,-6,-148,9,-4,11,-21,7,-34,-40,-64,-4,1,-9,-8,0,-52,-8,-18,-51,-41,-27,5,-31,4,-32,0,-60,-399,-27,-9,8,-28,0,-23,6,1,1,-16,36,-10,23,-65,1,-13,-10,-15,-72,-1,0,-7,-49,-5,-4,14,-11,-1,-2,-8,-17,8,10,-1,-40,-6,-74,-35,-2,-9,-6,-84,-15,-10,1,-8,7,4,-176,-1,-242,11,-1,2,-3,0,9,-160,-18,-113,-15,-43,-9,-16,-11,3,-39,2,-73,-47,6,-2,0,-7,-23,-11,-4,3,3,-3,0,11,-6,-37,-6,-574,-27,14,1,1,-44,-1,-21,-4,-14,-209,-48,0,25,-28,-36,-5,24,-3,-146,14,-481,-23,0,1,1,-4,-24,2,-1},
{-8,-12,-7,-10,-13,-4,1,-59,-16,-1,0,2,-30,-5,-451,-38,-3,-3,-15,1,-4,0,-5,-23,-7,-134,-9,0,-8,-9,-3,-26,-7,-5,-15,-71,-61,-164,-10,-13,-10,-1,-10,-44,-11,-8,-11,2,-2,-1,-12,-11,-74,0,-10,-7,-11,1,-2,-4,-1,-11,-10,-50,-79,-61,-4,-14,-11,-16,-16,-5,-8,-4,-5,-10,-25,-12,-3,0,5,-82,-2,-28,-55,-3,-6,2,-12,-14,-47,-7,-30,-9,-12,-12,-11,-7,-8,-15,1,-27,-29,-13,3,-3,-14,-3,-190,-12,3,5,-3,-21,2,-129,-7,1,-11,-44,-1,-6,-11,-10,1,2,-9,-11,-9,-5,0,-56,-9,-5,-17,-14,-8,-4,-7,4,-6,-6,-6,-3,-6,-4,-11,1,-29,-24,-14,0,0,-196,-1,-6,-14,-16,-8,-30,-12,7,-3,-2,-66,-9,2,-11,-6,-12,-25,-23,-4,6,-6,-9,-6,0,-6,-2,-4,-38,5,-10,-125,2,2,-11,-6,-20,-14,-34,-11,-6,-7,-5,-14,-29,-5,-8}
};

 NN  #(
    .output_number(output_number), 
    .input_number(input_number), 
    .width(width)) U_layer3(
    .clk(clk), 
    .rst_n(rst_n), 
    .enable(enable),
    .input_node(input_node),
    .bias(bias),
    .weight(weight), 
    .sum(internode), 
    .finish(finish)
);


relu #(
    .input_number(output_number),  
    .width(width)
    )U_relu4(
    .input_node(internode) , 
    .output_node(output_node)
    );



endmodule
